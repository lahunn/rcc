module rcc_vcore_clk_ctrl (
    output wire sys_clk,
    output wire sys_clk_pre,
    // signals connected to PAD 
    output      mco1,
    output      mco2,
    input       pad_rcc_eth_mii_tx_clk,
    input       pad_rcc_eth_mii_rx_clk,
    input       USB_PHY1,
    // signals connected to PWR 
    input       d3_deepsleep,
    output      c2_per_alloc_d1,
    output      c1_per_alloc_d2,
    // signals connected to CPU 
    input       c2_sleep,
    input       c2_deepsleep,
    input       c1_sleep,
    input       c1_deepsleep,
    output      rcc_c2_clk,
    output      rcc_fclk_c2,
    output      rcc_c2_systick_clk,
    output      rcc_c1_clk,
    output      rcc_fclk_c1,
    output      rcc_c1_systick_clk,
    // timer clocks
    output wire rcc_timx_ker_clk,
    output wire rcc_timy_ker_clk,
    output wire rcc_hrtimer_prescalar_clk,
    output wire sys_d1cpre_clk,
    output wire sys_hpre_clk,
    //rtc clocks
    output wire hse_rtc_clk,

    // stop mode signals
    input wire rcc_d1_stop,
    input wire rcc_d2_stop,
    input wire rcc_sys_stop,
    // signals connected to HSE
    input      hse_css_fail,
    input      hse_clk_pre,
    // lse lsi clock
    input      lse_clk,
    input      lsi_clk,
    // signals connected to HSI48 
    input      hsi48_clk,
    // signals connected to CSI
    input      csi_clk_pre,
    // signals connected to HSI
    input      hsi_origin_clk,

    // reset signals 
    input wire sys_rst_n,

    //bus clock signals
    output wire       rcc_axibridge_d1_clk,
    output wire       rcc_ahb3bridge_d1_clk,
    output wire       rcc_apb3bridge_d1_clk,
    output wire       rcc_ahb1bridge_d2_clk,
    output wire       rcc_ahb2bridge_d2_clk,
    output wire       rcc_apb1bridge_d2_clk,
    output wire       rcc_apb2bridge_d2_clk,
    output wire       rcc_ahb4bridge_d3_clk,
    output wire       rcc_apb4bridge_d3_clk,
    //pll , oscilator and pad clocks
    input  wire [1:0] pll_src_sel,
    input  wire       pll1_q_clk,
    input  wire       pll1_p_clk,
    input  wire       pll2_p_clk,
    input  wire       pll2_q_clk,
    input  wire       pll2_r_clk,
    input  wire       pll3_p_clk,
    input  wire       pll3_q_clk,
    input  wire       pll3_r_clk,
    input  wire       I2S_clk_IN,
    output            pll1_src_clk,
    output            pll2_src_clk,
    output            pll3_src_clk,

    //periperal enable signals
    input wire       rcc_c2_flash_en,
    input wire       rcc_c1_flash_lpen,
    input wire       rcc_c2_flash_lpen,
    input wire       rcc_c1_qspi_en,
    input wire       rcc_c2_qspi_en,
    input wire       rcc_c1_qspi_lpen,
    input wire       rcc_c2_qspi_lpen,
    input wire       rcc_c2_axisram_en,
    input wire       rcc_c1_axisram_lpen,
    input wire       rcc_c2_axisram_lpen,
    input wire       rcc_c1_fmc_en,
    input wire       rcc_c2_fmc_en,
    input wire       rcc_c1_fmc_lpen,
    input wire       rcc_c2_fmc_lpen,
    input wire       rcc_c1_dma2d_en,
    input wire       rcc_c2_dma2d_en,
    input wire       rcc_c1_dma2d_lpen,
    input wire       rcc_c2_dma2d_lpen,
    input wire       rcc_c1_mdma_en,
    input wire       rcc_c2_mdma_en,
    input wire       rcc_c1_mdma_lpen,
    input wire       rcc_c2_mdma_lpen,
    input wire       rcc_c1_ltdc_en,
    input wire       rcc_c2_ltdc_en,
    input wire       rcc_c1_ltdc_lpen,
    input wire       rcc_c2_ltdc_lpen,
    input wire       rcc_c2_itcm_en,
    input wire       rcc_c1_itcm_lpen,
    input wire       rcc_c2_itcm_lpen,
    input wire       rcc_c2_dtcm2_en,
    input wire       rcc_c1_dtcm2_lpen,
    input wire       rcc_c2_dtcm2_lpen,
    input wire       rcc_c2_dtcm1_en,
    input wire       rcc_c1_dtcm1_lpen,
    input wire       rcc_c2_dtcm1_lpen,
    input wire       rcc_c1_jpgdec_en,
    input wire       rcc_c2_jpgdec_en,
    input wire       rcc_c1_jpgdec_lpen,
    input wire       rcc_c2_jpgdec_lpen,
    input wire       rcc_c1_sdmmc1_en,
    input wire       rcc_c2_sdmmc1_en,
    input wire       rcc_c1_sdmmc1_lpen,
    input wire       rcc_c2_sdmmc1_lpen,
    input wire       rcc_c1_wwdg1_en,
    input wire       rcc_c2_wwdg1_en,
    input wire       rcc_c1_wwdg1_lpen,
    input wire       rcc_c2_wwdg1_lpen,
    input wire       rcc_c1_usb2ulpi_en,
    input wire       rcc_c2_usb2ulpi_en,
    input wire       rcc_c1_usb2ulpi_lpen,
    input wire       rcc_c2_usb2ulpi_lpen,
    input wire       rcc_c1_usb2otg_en,
    input wire       rcc_c2_usb2otg_en,
    input wire       rcc_c1_usb2otg_lpen,
    input wire       rcc_c2_usb2otg_lpen,
    input wire       rcc_c1_usb1ulpi_en,
    input wire       rcc_c2_usb1ulpi_en,
    input wire       rcc_c1_usb1ulpi_lpen,
    input wire       rcc_c2_usb1ulpi_lpen,
    input wire       rcc_c1_usb1otg_en,
    input wire       rcc_c2_usb1otg_en,
    input wire       rcc_c1_usb1otg_lpen,
    input wire       rcc_c2_usb1otg_lpen,
    input wire       rcc_c1_eth1rx_en,
    input wire       rcc_c2_eth1rx_en,
    input wire       rcc_c1_eth1rx_lpen,
    input wire       rcc_c2_eth1rx_lpen,
    input wire       rcc_c1_eth1tx_en,
    input wire       rcc_c2_eth1tx_en,
    input wire       rcc_c1_eth1tx_lpen,
    input wire       rcc_c2_eth1tx_lpen,
    input wire       rcc_c1_eth1mac_en,
    input wire       rcc_c2_eth1mac_en,
    input wire       rcc_c1_eth1mac_lpen,
    input wire       rcc_c2_eth1mac_lpen,
    input wire       rcc_c1_adc12_en,
    input wire       rcc_c2_adc12_en,
    input wire       rcc_c1_adc12_lpen,
    input wire       rcc_c2_adc12_lpen,
    input wire       rcc_c1_dma2_en,
    input wire       rcc_c2_dma2_en,
    input wire       rcc_c1_dma2_lpen,
    input wire       rcc_c2_dma2_lpen,
    input wire       rcc_c1_dma1_en,
    input wire       rcc_c2_dma1_en,
    input wire       rcc_c1_dma1_lpen,
    input wire       rcc_c2_dma1_lpen,
    input wire       rcc_c1_sram3_en,
    input wire       rcc_c1_sram3_lpen,
    input wire       rcc_c2_sram3_lpen,
    input wire       rcc_c1_sram2_en,
    input wire       rcc_c1_sram2_lpen,
    input wire       rcc_c2_sram2_lpen,
    input wire       rcc_c1_sram1_en,
    input wire       rcc_c1_sram1_lpen,
    input wire       rcc_c2_sram1_lpen,
    input wire       rcc_c1_sdmmc2_en,
    input wire       rcc_c2_sdmmc2_en,
    input wire       rcc_c1_sdmmc2_lpen,
    input wire       rcc_c2_sdmmc2_lpen,
    input wire       rcc_c1_rng_en,
    input wire       rcc_c2_rng_en,
    input wire       rcc_c1_rng_lpen,
    input wire       rcc_c2_rng_lpen,
    input wire       rcc_c1_hash_en,
    input wire       rcc_c2_hash_en,
    input wire       rcc_c1_hash_lpen,
    input wire       rcc_c2_hash_lpen,
    input wire       rcc_c1_crypt_en,
    input wire       rcc_c2_crypt_en,
    input wire       rcc_c1_crypt_lpen,
    input wire       rcc_c2_crypt_lpen,
    input wire       rcc_c1_dcmi_en,
    input wire       rcc_c2_dcmi_en,
    input wire       rcc_c1_dcmi_lpen,
    input wire       rcc_c2_dcmi_lpen,
    input wire       rcc_c1_uart8_en,
    input wire       rcc_c2_uart8_en,
    input wire       rcc_c1_uart8_lpen,
    input wire       rcc_c2_uart8_lpen,
    input wire       uart8_ker_clk_req,
    input wire       rcc_c1_uart7_en,
    input wire       rcc_c2_uart7_en,
    input wire       rcc_c1_uart7_lpen,
    input wire       rcc_c2_uart7_lpen,
    input wire       uart7_ker_clk_req,
    input wire       rcc_c1_dac12_en,
    input wire       rcc_c2_dac12_en,
    input wire       rcc_c1_dac12_lpen,
    input wire       rcc_c2_dac12_lpen,
    input wire       rcc_c1_hdmicec_en,
    input wire       rcc_c2_hdmicec_en,
    input wire       rcc_c1_hdmicec_lpen,
    input wire       rcc_c2_hdmicec_lpen,
    input wire       rcc_c1_i2c3_en,
    input wire       rcc_c2_i2c3_en,
    input wire       rcc_c1_i2c3_lpen,
    input wire       rcc_c2_i2c3_lpen,
    input wire       i2c3_ker_clk_req,
    input wire       rcc_c1_i2c2_en,
    input wire       rcc_c2_i2c2_en,
    input wire       rcc_c1_i2c2_lpen,
    input wire       rcc_c2_i2c2_lpen,
    input wire       i2c2_ker_clk_req,
    input wire       rcc_c1_i2c1_en,
    input wire       rcc_c2_i2c1_en,
    input wire       rcc_c1_i2c1_lpen,
    input wire       rcc_c2_i2c1_lpen,
    input wire       i2c1_ker_clk_req,
    input wire       rcc_c1_uart5_en,
    input wire       rcc_c2_uart5_en,
    input wire       rcc_c1_uart5_lpen,
    input wire       rcc_c2_uart5_lpen,
    input wire       uart5_ker_clk_req,
    input wire       rcc_c1_uart4_en,
    input wire       rcc_c2_uart4_en,
    input wire       rcc_c1_uart4_lpen,
    input wire       rcc_c2_uart4_lpen,
    input wire       uart4_ker_clk_req,
    input wire       rcc_c1_usart3_en,
    input wire       rcc_c2_usart3_en,
    input wire       rcc_c1_usart3_lpen,
    input wire       rcc_c2_usart3_lpen,
    input wire       usart3_ker_clk_req,
    input wire       rcc_c1_usart2_en,
    input wire       rcc_c2_usart2_en,
    input wire       rcc_c1_usart2_lpen,
    input wire       rcc_c2_usart2_lpen,
    input wire       usart2_ker_clk_req,
    input wire       rcc_c1_spdifrx_en,
    input wire       rcc_c2_spdifrx_en,
    input wire       rcc_c1_spdifrx_lpen,
    input wire       rcc_c2_spdifrx_lpen,
    input wire       rcc_c1_spi3_en,
    input wire       rcc_c2_spi3_en,
    input wire       rcc_c1_spi3_lpen,
    input wire       rcc_c2_spi3_lpen,
    input wire       rcc_c1_spi2_en,
    input wire       rcc_c2_spi2_en,
    input wire       rcc_c1_spi2_lpen,
    input wire       rcc_c2_spi2_lpen,
    input wire       rcc_c1_wwdg2_en,
    input wire       rcc_c2_wwdg2_en,
    input wire       rcc_c1_wwdg2_lpen,
    input wire       rcc_c2_wwdg2_lpen,
    input wire       rcc_c1_lptim1_en,
    input wire       rcc_c2_lptim1_en,
    input wire       rcc_c1_lptim1_lpen,
    input wire       rcc_c2_lptim1_lpen,
    input wire       rcc_c1_tim14_en,
    input wire       rcc_c2_tim14_en,
    input wire       rcc_c1_tim14_lpen,
    input wire       rcc_c2_tim14_lpen,
    input wire       rcc_c1_tim13_en,
    input wire       rcc_c2_tim13_en,
    input wire       rcc_c1_tim13_lpen,
    input wire       rcc_c2_tim13_lpen,
    input wire       rcc_c1_tim12_en,
    input wire       rcc_c2_tim12_en,
    input wire       rcc_c1_tim12_lpen,
    input wire       rcc_c2_tim12_lpen,
    input wire       rcc_c1_tim7_en,
    input wire       rcc_c2_tim7_en,
    input wire       rcc_c1_tim7_lpen,
    input wire       rcc_c2_tim7_lpen,
    input wire       rcc_c1_tim6_en,
    input wire       rcc_c2_tim6_en,
    input wire       rcc_c1_tim6_lpen,
    input wire       rcc_c2_tim6_lpen,
    input wire       rcc_c1_tim5_en,
    input wire       rcc_c2_tim5_en,
    input wire       rcc_c1_tim5_lpen,
    input wire       rcc_c2_tim5_lpen,
    input wire       rcc_c1_tim4_en,
    input wire       rcc_c2_tim4_en,
    input wire       rcc_c1_tim4_lpen,
    input wire       rcc_c2_tim4_lpen,
    input wire       rcc_c1_tim3_en,
    input wire       rcc_c2_tim3_en,
    input wire       rcc_c1_tim3_lpen,
    input wire       rcc_c2_tim3_lpen,
    input wire       rcc_c1_tim2_en,
    input wire       rcc_c2_tim2_en,
    input wire       rcc_c1_tim2_lpen,
    input wire       rcc_c2_tim2_lpen,
    input wire       rcc_c1_fdcan_en,
    input wire       rcc_c2_fdcan_en,
    input wire       rcc_c1_fdcan_lpen,
    input wire       rcc_c2_fdcan_lpen,
    input wire       rcc_c1_mdios_en,
    input wire       rcc_c2_mdios_en,
    input wire       rcc_c1_mdios_lpen,
    input wire       rcc_c2_mdios_lpen,
    input wire       rcc_c1_opamp_en,
    input wire       rcc_c2_opamp_en,
    input wire       rcc_c1_opamp_lpen,
    input wire       rcc_c2_opamp_lpen,
    input wire       rcc_c1_swpmi_en,
    input wire       rcc_c2_swpmi_en,
    input wire       rcc_c1_swpmi_lpen,
    input wire       rcc_c2_swpmi_lpen,
    input wire       rcc_c1_crs_en,
    input wire       rcc_c2_crs_en,
    input wire       rcc_c1_crs_lpen,
    input wire       rcc_c2_crs_lpen,
    input wire       rcc_c1_hrtim_en,
    input wire       rcc_c2_hrtim_en,
    input wire       rcc_c1_hrtim_lpen,
    input wire       rcc_c2_hrtim_lpen,
    input wire       rcc_c1_dfsdm1_en,
    input wire       rcc_c2_dfsdm1_en,
    input wire       rcc_c1_dfsdm1_lpen,
    input wire       rcc_c2_dfsdm1_lpen,
    input wire       rcc_c1_sai3_en,
    input wire       rcc_c2_sai3_en,
    input wire       rcc_c1_sai3_lpen,
    input wire       rcc_c2_sai3_lpen,
    input wire       rcc_c1_sai2_en,
    input wire       rcc_c2_sai2_en,
    input wire       rcc_c1_sai2_lpen,
    input wire       rcc_c2_sai2_lpen,
    input wire       rcc_c1_sai1_en,
    input wire       rcc_c2_sai1_en,
    input wire       rcc_c1_sai1_lpen,
    input wire       rcc_c2_sai1_lpen,
    input wire       rcc_c1_spi5_en,
    input wire       rcc_c2_spi5_en,
    input wire       rcc_c1_spi5_lpen,
    input wire       rcc_c2_spi5_lpen,
    input wire       rcc_c1_tim17_en,
    input wire       rcc_c2_tim17_en,
    input wire       rcc_c1_tim17_lpen,
    input wire       rcc_c2_tim17_lpen,
    input wire       rcc_c1_tim16_en,
    input wire       rcc_c2_tim16_en,
    input wire       rcc_c1_tim16_lpen,
    input wire       rcc_c2_tim16_lpen,
    input wire       rcc_c1_tim15_en,
    input wire       rcc_c2_tim15_en,
    input wire       rcc_c1_tim15_lpen,
    input wire       rcc_c2_tim15_lpen,
    input wire       rcc_c1_spi4_en,
    input wire       rcc_c2_spi4_en,
    input wire       rcc_c1_spi4_lpen,
    input wire       rcc_c2_spi4_lpen,
    input wire       rcc_c1_spi1_en,
    input wire       rcc_c2_spi1_en,
    input wire       rcc_c1_spi1_lpen,
    input wire       rcc_c2_spi1_lpen,
    input wire       rcc_c1_usart6_en,
    input wire       rcc_c2_usart6_en,
    input wire       rcc_c1_usart6_lpen,
    input wire       rcc_c2_usart6_lpen,
    input wire       usart6_ker_clk_req,
    input wire       rcc_c1_usart1_en,
    input wire       rcc_c2_usart1_en,
    input wire       rcc_c1_usart1_lpen,
    input wire       rcc_c2_usart1_lpen,
    input wire       usart1_ker_clk_req,
    input wire       rcc_c1_tim8_en,
    input wire       rcc_c2_tim8_en,
    input wire       rcc_c1_tim8_lpen,
    input wire       rcc_c2_tim8_lpen,
    input wire       rcc_c1_tim1_en,
    input wire       rcc_c2_tim1_en,
    input wire       rcc_c1_tim1_lpen,
    input wire       rcc_c2_tim1_lpen,
    input wire       rcc_c1_sram4_lpen,
    input wire       rcc_c2_sram4_lpen,
    input wire       rcc_sram4_amen,
    input wire       rcc_c1_bkpram_en,
    input wire       rcc_c2_bkpram_en,
    input wire       rcc_c1_bkpram_lpen,
    input wire       rcc_c2_bkpram_lpen,
    input wire       rcc_bkpram_amen,
    input wire       rcc_c1_hsem_en,
    input wire       rcc_c2_hsem_en,
    input wire       rcc_c1_adc3_en,
    input wire       rcc_c2_adc3_en,
    input wire       rcc_c1_adc3_lpen,
    input wire       rcc_c2_adc3_lpen,
    input wire       rcc_adc3_amen,
    input wire       rcc_c1_bdma_en,
    input wire       rcc_c2_bdma_en,
    input wire       rcc_c1_bdma_lpen,
    input wire       rcc_c2_bdma_lpen,
    input wire       rcc_bdma_amen,
    input wire       rcc_c1_crc_en,
    input wire       rcc_c2_crc_en,
    input wire       rcc_c1_crc_lpen,
    input wire       rcc_c2_crc_lpen,
    input wire       rcc_crc_amen,
    input wire       rcc_c1_gpiok_en,
    input wire       rcc_c2_gpiok_en,
    input wire       rcc_c1_gpiok_lpen,
    input wire       rcc_c2_gpiok_lpen,
    input wire       rcc_c1_gpioj_en,
    input wire       rcc_c2_gpioj_en,
    input wire       rcc_c1_gpioj_lpen,
    input wire       rcc_c2_gpioj_lpen,
    input wire       rcc_c1_gpioi_en,
    input wire       rcc_c2_gpioi_en,
    input wire       rcc_c1_gpioi_lpen,
    input wire       rcc_c2_gpioi_lpen,
    input wire       rcc_c1_gpioh_en,
    input wire       rcc_c2_gpioh_en,
    input wire       rcc_c1_gpioh_lpen,
    input wire       rcc_c2_gpioh_lpen,
    input wire       rcc_c1_gpiog_en,
    input wire       rcc_c2_gpiog_en,
    input wire       rcc_c1_gpiog_lpen,
    input wire       rcc_c2_gpiog_lpen,
    input wire       rcc_c1_gpiof_en,
    input wire       rcc_c2_gpiof_en,
    input wire       rcc_c1_gpiof_lpen,
    input wire       rcc_c2_gpiof_lpen,
    input wire       rcc_c1_gpioe_en,
    input wire       rcc_c2_gpioe_en,
    input wire       rcc_c1_gpioe_lpen,
    input wire       rcc_c2_gpioe_lpen,
    input wire       rcc_c1_gpiod_en,
    input wire       rcc_c2_gpiod_en,
    input wire       rcc_c1_gpiod_lpen,
    input wire       rcc_c2_gpiod_lpen,
    input wire       rcc_c1_gpioc_en,
    input wire       rcc_c2_gpioc_en,
    input wire       rcc_c1_gpioc_lpen,
    input wire       rcc_c2_gpioc_lpen,
    input wire       rcc_c1_gpiob_en,
    input wire       rcc_c2_gpiob_en,
    input wire       rcc_c1_gpiob_lpen,
    input wire       rcc_c2_gpiob_lpen,
    input wire       rcc_c1_gpioa_en,
    input wire       rcc_c2_gpioa_en,
    input wire       rcc_c1_gpioa_lpen,
    input wire       rcc_c2_gpioa_lpen,
    input wire       rcc_c1_sai4_en,
    input wire       rcc_c2_sai4_en,
    input wire       rcc_c1_sai4_lpen,
    input wire       rcc_c2_sai4_lpen,
    input wire       rcc_sai4_amen,
    input wire       rcc_c1_rtc_en,
    input wire       rcc_c2_rtc_en,
    input wire       rcc_c1_rtc_lpen,
    input wire       rcc_c2_rtc_lpen,
    input wire       rcc_rtc_amen,
    input wire       rcc_c1_vref_en,
    input wire       rcc_c2_vref_en,
    input wire       rcc_c1_vref_lpen,
    input wire       rcc_c2_vref_lpen,
    input wire       rcc_vref_amen,
    input wire       rcc_c1_comp12_en,
    input wire       rcc_c2_comp12_en,
    input wire       rcc_c1_comp12_lpen,
    input wire       rcc_c2_comp12_lpen,
    input wire       rcc_comp12_amen,
    input wire       rcc_c1_lptim5_en,
    input wire       rcc_c2_lptim5_en,
    input wire       rcc_c1_lptim5_lpen,
    input wire       rcc_c2_lptim5_lpen,
    input wire       rcc_lptim5_amen,
    input wire       rcc_c1_lptim4_en,
    input wire       rcc_c2_lptim4_en,
    input wire       rcc_c1_lptim4_lpen,
    input wire       rcc_c2_lptim4_lpen,
    input wire       rcc_lptim4_amen,
    input wire       rcc_c1_lptim3_en,
    input wire       rcc_c2_lptim3_en,
    input wire       rcc_c1_lptim3_lpen,
    input wire       rcc_c2_lptim3_lpen,
    input wire       rcc_lptim3_amen,
    input wire       rcc_c1_lptim2_en,
    input wire       rcc_c2_lptim2_en,
    input wire       rcc_c1_lptim2_lpen,
    input wire       rcc_c2_lptim2_lpen,
    input wire       rcc_lptim2_amen,
    input wire       rcc_c1_i2c4_en,
    input wire       rcc_c2_i2c4_en,
    input wire       rcc_c1_i2c4_lpen,
    input wire       rcc_c2_i2c4_lpen,
    input wire       rcc_i2c4_amen,
    input wire       i2c4_ker_clk_req,
    input wire       rcc_c1_spi6_en,
    input wire       rcc_c2_spi6_en,
    input wire       rcc_c1_spi6_lpen,
    input wire       rcc_c2_spi6_lpen,
    input wire       rcc_spi6_amen,
    input wire       rcc_c1_lpuart1_en,
    input wire       rcc_c2_lpuart1_en,
    input wire       rcc_c1_lpuart1_lpen,
    input wire       rcc_c2_lpuart1_lpen,
    input wire       rcc_lpuart1_amen,
    input wire       lpuart1_ker_clk_req,
    input wire       rcc_c1_syscfg_en,
    input wire       rcc_c2_syscfg_en,
    input wire       rcc_c1_syscfg_lpen,
    input wire       rcc_c2_syscfg_lpen,
    //clk sel signals from register
    input wire [1:0] qspisel,
    input wire [1:0] fmcsel,
    input wire       sdmmcsel,
    input wire [1:0] usbsel,
    input wire [1:0] adcsel,
    input wire [1:0] rngsel,
    input wire [1:0] cecsel,
    input wire [1:0] i2c123sel,
    input wire [2:0] usart234578sel,
    input wire [1:0] spdifsel,
    input wire [2:0] lptim1sel,
    input wire [1:0] fdcansel,
    input wire       swpmisel,
    input wire [2:0] sai1sel,
    input wire       dfsdm1sel,
    input wire [2:0] sai23sel,
    input wire [2:0] spi45sel,
    input wire [2:0] spi123sel,
    input wire [2:0] usart16sel,
    input wire [2:0] sai4asel,
    input wire [2:0] sai4bsel,
    input wire [2:0] lptim345sel,
    input wire [2:0] lptim2sel,
    input wire [1:0] i2c4sel,
    input wire [2:0] spi6sel,
    input wire [2:0] lpuart1sel,




    // per_ker_clk_control Outputs
    //per_ker_clk_control region
    output wire rcc_rtc_pclk,
    output wire rcc_flash_aclk,
    output wire rcc_flash_hclk,
    output wire rcc_qspi_aclk,
    output wire rcc_qspi_hclk,
    output wire rcc_qspi_ker_clk,
    output wire rcc_axisram_aclk,
    output wire rcc_fmc_aclk,
    output wire rcc_fmc_hclk,
    output wire rcc_fmc_ker_clk,
    output wire rcc_dma2d_aclk,
    output wire rcc_dma2d_hclk,
    output wire rcc_mdma_aclk,
    output wire rcc_mdma_hclk,
    output wire rcc_ltdc_aclk,
    output wire rcc_ltdc_pclk,
    output wire rcc_ltdc_ker_clk,
    output wire rcc_ramecc1_hclk,
    output wire rcc_gpv_hclk,
    output wire rcc_itcm_hclk,
    output wire rcc_dtcm2_hclk,
    output wire rcc_dtcm1_hclk,
    output wire rcc_jpgdec_hclk,
    output wire rcc_sdmmc1_hclk,
    output wire rcc_sdmmc1_ker_clk,
    output wire rcc_wwdg1_pclk,
    output wire rcc_usb2ulpi_hclk,
    output wire rcc_usb2otg_hclk,
    output wire rcc_usb2otg_ker_clk,
    output wire rcc_usb1ulpi_hclk,
    output wire rcc_usb1ulpi_ker_clk,
    output wire rcc_usb1otg_hclk,
    output wire rcc_usb1otg_ker_clk,
    output wire rcc_eth1rx_hclk,
    output wire rcc_eth1tx_hclk,
    output wire rcc_eth1mac_hclk,
    output wire rcc_adc12_hclk,
    output wire rcc_adc12_ker_clk,
    output wire rcc_dma2_hclk,
    output wire rcc_dma1_hclk,
    output wire rcc_sram3_hclk,
    output wire rcc_sram2_hclk,
    output wire rcc_sram1_hclk,
    output wire rcc_sdmmc2_hclk,
    output wire rcc_sdmmc2_ker_clk,
    output wire rcc_rng_hclk,
    output wire rcc_rng_ker_clk,
    output wire rcc_hash_hclk,
    output wire rcc_crypt_hclk,
    output wire rcc_dcmi_hclk,
    output wire rcc_ramecc2_hclk,
    output wire rcc_uart8_pclk,
    output wire rcc_uart8_ker_clk,
    output wire rcc_uart7_pclk,
    output wire rcc_uart7_ker_clk,
    output wire rcc_dac12_pclk,
    output wire rcc_hdmicec_pclk,
    output wire rcc_hdmicec_ker_clk,
    output wire rcc_i2c3_pclk,
    output wire rcc_i2c3_ker_clk,
    output wire rcc_i2c2_pclk,
    output wire rcc_i2c2_ker_clk,
    output wire rcc_i2c1_pclk,
    output wire rcc_i2c1_ker_clk,
    output wire rcc_uart5_pclk,
    output wire rcc_uart5_ker_clk,
    output wire rcc_uart4_pclk,
    output wire rcc_uart4_ker_clk,
    output wire rcc_usart3_pclk,
    output wire rcc_usart3_ker_clk,
    output wire rcc_usart2_pclk,
    output wire rcc_usart2_ker_clk,
    output wire rcc_spdifrx_pclk,
    output wire rcc_spdifrx_ker_clk,
    output wire rcc_spi3_pclk,
    output wire rcc_spi3_ker_clk,
    output wire rcc_spi2_pclk,
    output wire rcc_spi2_ker_clk,
    output wire rcc_wwdg2_pclk,
    output wire rcc_lptim1_pclk,
    output wire rcc_lptim1_ker_clk,
    output wire rcc_tim14_pclk,
    output wire rcc_tim14_ker_clk,
    output wire rcc_tim13_pclk,
    output wire rcc_tim13_ker_clk,
    output wire rcc_tim12_pclk,
    output wire rcc_tim12_ker_clk,
    output wire rcc_tim7_pclk,
    output wire rcc_tim7_ker_clk,
    output wire rcc_tim6_pclk,
    output wire rcc_tim6_ker_clk,
    output wire rcc_tim5_pclk,
    output wire rcc_tim5_ker_clk,
    output wire rcc_tim4_pclk,
    output wire rcc_tim4_ker_clk,
    output wire rcc_tim3_pclk,
    output wire rcc_tim3_ker_clk,
    output wire rcc_tim2_pclk,
    output wire rcc_tim2_ker_clk,
    output wire rcc_fdcan_pclk,
    output wire rcc_fdcan_ker_clk,
    output wire rcc_mdios_pclk,
    output wire rcc_opamp_pclk,
    output wire rcc_swpmi_pclk,
    output wire rcc_swpmi_ker_clk,
    output wire rcc_crs_pclk,
    output wire rcc_hrtim_pclk,
    output wire rcc_hrtim_ker_clk,
    output wire rcc_dfsdm1_pclk,
    output wire rcc_dfsdm1_ker_clk_0,
    output wire rcc_dfsdm1_ker_clk_1,
    output wire rcc_sai3_pclk,
    output wire rcc_sai3_ker_clk,
    output wire rcc_sai2_pclk,
    output wire rcc_sai2_ker_clk,
    output wire rcc_sai1_pclk,
    output wire rcc_sai1_ker_clk,
    output wire rcc_spi5_pclk,
    output wire rcc_spi5_ker_clk,
    output wire rcc_tim17_pclk,
    output wire rcc_tim17_ker_clk,
    output wire rcc_tim16_pclk,
    output wire rcc_tim16_ker_clk,
    output wire rcc_tim15_pclk,
    output wire rcc_tim15_ker_clk,
    output wire rcc_spi4_pclk,
    output wire rcc_spi4_ker_clk,
    output wire rcc_spi1_pclk,
    output wire rcc_spi1_ker_clk,
    output wire rcc_usart6_pclk,
    output wire rcc_usart6_ker_clk,
    output wire rcc_usart1_pclk,
    output wire rcc_usart1_ker_clk,
    output wire rcc_tim8_pclk,
    output wire rcc_tim8_ker_clk,
    output wire rcc_tim1_pclk,
    output wire rcc_tim1_ker_clk,
    output wire rcc_sram4_hclk,
    output wire rcc_bkpram_hclk,
    output wire rcc_ramecc3_hclk,
    output wire rcc_hsem_hclk,
    output wire rcc_adc3_hclk,
    output wire rcc_adc3_ker_clk,
    output wire rcc_bdma_hclk,
    output wire rcc_crc_hclk,
    output wire rcc_gpiok_hclk,
    output wire rcc_gpioj_hclk,
    output wire rcc_gpioi_hclk,
    output wire rcc_gpioh_hclk,
    output wire rcc_gpiog_hclk,
    output wire rcc_gpiof_hclk,
    output wire rcc_gpioe_hclk,
    output wire rcc_gpiod_hclk,
    output wire rcc_gpioc_hclk,
    output wire rcc_gpiob_hclk,
    output wire rcc_gpioa_hclk,
    output wire rcc_rcc_hclk,
    output wire rcc_pwr_hclk,
    output wire rcc_sai4_pclk,
    output wire rcc_sai4_ker_clk_0,
    output wire rcc_sai4_ker_clk_1,
    output wire rcc_vref_pclk,
    output wire rcc_comp12_pclk,
    output wire rcc_lptim5_pclk,
    output wire rcc_lptim5_ker_clk,
    output wire rcc_lptim4_pclk,
    output wire rcc_lptim4_ker_clk,
    output wire rcc_lptim3_pclk,
    output wire rcc_lptim3_ker_clk,
    output wire rcc_lptim2_pclk,
    output wire rcc_lptim2_ker_clk,
    output wire rcc_i2c4_pclk,
    output wire rcc_i2c4_ker_clk,
    output wire rcc_spi6_pclk,
    output wire rcc_spi6_ker_clk,
    output wire rcc_lpuart1_pclk,
    output wire rcc_lpuart1_ker_clk,
    output wire rcc_syscfg_pclk,
    output wire rcc_iwdg2_pclk,
    output wire rcc_iwdg1_pclk,
    output wire rcc_exti_pclk,
    //end per_ker_clk_control region

    //rcc_sys_async_reset_clk_gate enable signals
    input        d1_clk_arcg_en,
    input        d2_clk_arcg_en,
    input        cpu1_clk_arcg_en,
    input        cpu2_clk_arcg_en,
    input        sys_clk_arcg_en,
    input        rcc_flash_arcg_clk_en,
    input        rcc_qspi_arcg_clk_en,
    input        rcc_axisram_arcg_clk_en,
    input        rcc_fmc_arcg_clk_en,
    input        rcc_dma2d_arcg_clk_en,
    input        rcc_mdma_arcg_clk_en,
    input        rcc_ltdc_arcg_clk_en,
    input        rcc_ramecc1_arcg_clk_en,
    input        rcc_gpv_arcg_clk_en,
    input        rcc_itcm_arcg_clk_en,
    input        rcc_dtcm2_arcg_clk_en,
    input        rcc_dtcm1_arcg_clk_en,
    input        rcc_jpgdec_arcg_clk_en,
    input        rcc_sdmmc1_arcg_clk_en,
    input        rcc_wwdg1_arcg_clk_en,
    input        rcc_usb2ulpi_arcg_clk_en,
    input        rcc_usb2otg_arcg_clk_en,
    input        rcc_usb1ulpi_arcg_clk_en,
    input        rcc_usb1otg_arcg_clk_en,
    input        rcc_eth1rx_arcg_clk_en,
    input        rcc_eth1tx_arcg_clk_en,
    input        rcc_eth1mac_arcg_clk_en,
    input        rcc_adc12_arcg_clk_en,
    input        rcc_dma2_arcg_clk_en,
    input        rcc_dma1_arcg_clk_en,
    input        rcc_sram3_arcg_clk_en,
    input        rcc_sram2_arcg_clk_en,
    input        rcc_sram1_arcg_clk_en,
    input        rcc_sdmmc2_arcg_clk_en,
    input        rcc_rng_arcg_clk_en,
    input        rcc_hash_arcg_clk_en,
    input        rcc_crypt_arcg_clk_en,
    input        rcc_dcmi_arcg_clk_en,
    input        rcc_ramecc2_arcg_clk_en,
    input        rcc_uart8_arcg_clk_en,
    input        rcc_uart7_arcg_clk_en,
    input        rcc_dac12_arcg_clk_en,
    input        rcc_hdmicec_arcg_clk_en,
    input        rcc_i2c3_arcg_clk_en,
    input        rcc_i2c2_arcg_clk_en,
    input        rcc_i2c1_arcg_clk_en,
    input        rcc_uart5_arcg_clk_en,
    input        rcc_uart4_arcg_clk_en,
    input        rcc_usart3_arcg_clk_en,
    input        rcc_usart2_arcg_clk_en,
    input        rcc_spdifrx_arcg_clk_en,
    input        rcc_spi3_arcg_clk_en,
    input        rcc_spi2_arcg_clk_en,
    input        rcc_wwdg2_arcg_clk_en,
    input        rcc_lptim1_arcg_clk_en,
    input        rcc_tim14_arcg_clk_en,
    input        rcc_tim13_arcg_clk_en,
    input        rcc_tim12_arcg_clk_en,
    input        rcc_tim7_arcg_clk_en,
    input        rcc_tim6_arcg_clk_en,
    input        rcc_tim5_arcg_clk_en,
    input        rcc_tim4_arcg_clk_en,
    input        rcc_tim3_arcg_clk_en,
    input        rcc_tim2_arcg_clk_en,
    input        rcc_fdcan_arcg_clk_en,
    input        rcc_mdios_arcg_clk_en,
    input        rcc_opamp_arcg_clk_en,
    input        rcc_swpmi_arcg_clk_en,
    input        rcc_crs_arcg_clk_en,
    input        rcc_hrtim_arcg_clk_en,
    input        rcc_dfsdm1_arcg_clk_en,
    input        rcc_sai3_arcg_clk_en,
    input        rcc_sai2_arcg_clk_en,
    input        rcc_sai1_arcg_clk_en,
    input        rcc_spi5_arcg_clk_en,
    input        rcc_tim17_arcg_clk_en,
    input        rcc_tim16_arcg_clk_en,
    input        rcc_tim15_arcg_clk_en,
    input        rcc_spi4_arcg_clk_en,
    input        rcc_spi1_arcg_clk_en,
    input        rcc_usart6_arcg_clk_en,
    input        rcc_usart1_arcg_clk_en,
    input        rcc_tim8_arcg_clk_en,
    input        rcc_tim1_arcg_clk_en,
    input        rcc_sram4_arcg_clk_en,
    input        rcc_bkpram_arcg_clk_en,
    input        rcc_ramecc3_arcg_clk_en,
    input        rcc_hsem_arcg_clk_en,
    input        rcc_adc3_arcg_clk_en,
    input        rcc_bdma_arcg_clk_en,
    input        rcc_crc_arcg_clk_en,
    input        rcc_gpiok_arcg_clk_en,
    input        rcc_gpioj_arcg_clk_en,
    input        rcc_gpioi_arcg_clk_en,
    input        rcc_gpioh_arcg_clk_en,
    input        rcc_gpiog_arcg_clk_en,
    input        rcc_gpiof_arcg_clk_en,
    input        rcc_gpioe_arcg_clk_en,
    input        rcc_gpiod_arcg_clk_en,
    input        rcc_gpioc_arcg_clk_en,
    input        rcc_gpiob_arcg_clk_en,
    input        rcc_gpioa_arcg_clk_en,
    input        rcc_rcc_arcg_clk_en,
    input        rcc_pwr_arcg_clk_en,
    input        rcc_sai4_arcg_clk_en,
    input        rcc_rtc_arcg_clk_en,
    input        rcc_vref_arcg_clk_en,
    input        rcc_comp12_arcg_clk_en,
    input        rcc_lptim5_arcg_clk_en,
    input        rcc_lptim4_arcg_clk_en,
    input        rcc_lptim3_arcg_clk_en,
    input        rcc_lptim2_arcg_clk_en,
    input        rcc_i2c4_arcg_clk_en,
    input        rcc_spi6_arcg_clk_en,
    input        rcc_lpuart1_arcg_clk_en,
    input        rcc_syscfg_arcg_clk_en,
    input        rcc_iwdg2_arcg_clk_en,
    input        rcc_iwdg1_arcg_clk_en,
    input        rcc_exti_arcg_clk_en,
    //end rcc_sys_async_reset_clk_gate region
    //signals from eth and to eth
    input        eth_rcc_fes,
    input        eth_rcc_epis_2,
    output       rcc_eth_mii_tx_clk,
    output       rcc_eth_mii_rx_clk,
    output       rcc_eth_rmii_ref_clk,
    // register signals
    input  [2:0] mco1sel,
    input  [2:0] mco2sel,
    input  [3:0] mco1pre,
    input  [3:0] mco2pre,
    input  [5:0] rtcpre,
    input  [1:0] hsidiv,
    input  [1:0] sys_clk_sw,
    input  [3:0] d1cpre,
    input  [2:0] d1ppre,
    input  [3:0] hpre,
    input  [2:0] d2ppre1,
    input  [2:0] d2ppre2,
    input  [2:0] d3ppre,
    input        timpre,
    input        hrtimsel,
    input  [1:0] clkpersel,
    input  [5:0] divm1,
    input  [5:0] divm2,
    input  [5:0] divm3
);


  //////////////////////////////////
  //signals definition
  //////////////////////////////////
  wire hse_clk_en;
  wire hse_clk;

  wire hsi_clk_pre;  // hsi_clk is the clock before gate
  wire hsi_clk;
  wire hsi_ker_clk;
  wire hsi_clk_en;
  wire hsi_ker_clk_en;

  wire csi_clk;
  wire csi_clk_en;
  wire csi_ker_clk;
  wire csi_ker_clk_en;

  wire per_clk;

  wire pll_src_clk;

  wire hsi_ker_clk_req;
  wire csi_ker_clk_req;

  wire mco1_clk_pre;
  wire mco2_clk_pre;

  //////////////////////////////////
  // 

  //////////////////////////////////
  // HSI CSI clock control /////////
  //////////////////////////////////

  assign hsi_clk_en     = ~rcc_sys_stop;
  assign hsi_ker_clk_en = ~rcc_sys_stop | hsi_ker_clk_req;
  assign csi_clk_en     = ~rcc_sys_stop;
  assign csi_ker_clk_en = csi_clk_en | csi_ker_clk_req;


  assign hse_clk_en     = ~hse_css_fail;

  //////////////////////////////////
  // MCO clock out
  //////////////////////////////////

  mux_N_to_1 #(
      .N(5),
      .m(3)
  ) mco1_clk_switch_cell (
      .inp   ({hsi48_clk, pll1_q_clk, hse_clk, lse_clk, hsi_clk}),
      .select(mco1sel),

      .out(mco1_clk_pre)
  );

  div_odd_even #(
      .MAX_DIV_FAC(15)
  ) mco1_clk_divider (
      .clk_in (mco1_clk_pre),
      .rst_n  (sys_rst_n),
      .div_sel(mco1pre),

      .clk_out(mco1)
  );

  mux_N_to_1 #(
      .N(6),
      .m(3)
  ) mco2_clk_switch_cell (
      .inp   ({lsi_clk, csi_clk, pll1_p_clk, hse_clk, pll2_p_clk, sys_clk}),
      .select(mco2sel),

      .out(mco2_clk_pre)
  );

  div_odd_even #(
      .MAX_DIV_FAC(15)
  ) mco2_clk_divider (
      .clk_in (mco2_clk_pre),
      .rst_n  (sys_rst_n),
      .div_sel(mco2pre),

      .clk_out(mco2)
  );


  //////////////////////////////////
  // hse_rtc_clk generate
  //////////////////////////////////

  div_odd_even #(
      .MAX_DIV_FAC(63)
  ) hse_rtc_clk_div (
      .clk_in (hse_clk_pre),
      .rst_n  (sys_rst_n),
      .div_sel(rtcpre),

      .clk_out(hse_rtc_clk)
  );


  //////////////////////////////////
  // hsi_div
  //////////////////////////////////

  div_x_stage #(
      .STAGE_NUM      (3),
      .IS_STAGE_REMOVE(0),
      .STAGE_REMOVED  (0)
  ) hsi_clk_div (
      .clk_in (hsi_origin_clk),
      .rst_n  (sys_rst_n),
      .div_sel(hsidiv),

      .clk_out(hsi_clk_pre)
  );

  ////////////////////////////////
  //hsi clk gate
  ///////////////////////////////

  rcc_clk_gate_cell hsi_clk_gate (
      .clk_in(hsi_clk_pre),
      .clk_en(hsi_clk_en),

      .clk_out(hsi_clk)
  );

  rcc_clk_gate_cell hsi_ker_clk_gate (
      .clk_in(hsi_clk_pre),
      .clk_en(hsi_ker_clk_en),

      .clk_out(hsi_ker_clk)
  );

  //////////////////////////////
  //hse clk gate
  /////////////////////////////
  rcc_clk_gate_cell hse_clk_gate (
      .clk_in (hse_clk_pre),
      .clk_en (hse_clk_en),
      .clk_out(hse_clk)
  );

  ////////////////////////////
  //csi clock gate
  ///////////////////////////

  rcc_clk_gate_cell csi_clk_gate (
      .clk_in(csi_clk_pre),
      .clk_en(csi_clk_en),

      .clk_out(csi_clk)
  );

  rcc_clk_gate_cell csi_ker_clk_gate (
      .clk_in(csi_clk_pre),
      .clk_en(csi_ker_clk_en),

      .clk_out(csi_ker_clk)
  );

  ////////////////////////////
  //per_clk selection
  ///////////////////////////
  glitch_free_clk_switch #(
      .CLK_NUM(3)
  ) per_clk_switch (
      .clk_in ({hse_clk, csi_ker_clk, hsi_ker_clk}),
      .rst_n  (sys_rst_n),
      .sel    (clkpersel),
      .clk_out(per_clk)
  );



  ////////////////////////////
  //pll source clock generate
  ///////////////////////////

  glitch_free_clk_switch #(
      .CLK_NUM(3)
  ) pll_src_clk_switch (
      .clk_in({hse_clk, csi_clk, hsi_clk}),
      .rst_n (sys_rst_n),
      .sel   (pll_src_sel),

      .clk_out(pll_src_clk)
  );

  div_odd_even #(
      .MAX_DIV_FAC(63)
  ) pll1_src_clk_div (
      .clk_in (pll_src_clk),
      .rst_n  (sys_rst_n),
      .div_sel(divm1),

      .clk_out(pll1_src_clk)
  );

  div_odd_even #(
      .MAX_DIV_FAC(63)
  ) pll2_src_clk_div (
      .clk_in (pll_src_clk),
      .rst_n  (sys_rst_n),
      .div_sel(divm2),

      .clk_out(pll2_src_clk)
  );

  div_odd_even #(
      .MAX_DIV_FAC(63)
  ) pll3_src_clk_div (
      .clk_in (pll_src_clk),
      .rst_n  (sys_rst_n),
      .div_sel(divm3),

      .clk_out(pll3_src_clk)
  );

  rcc_sys_clk_gen u_rcc_sys_clk_gen (
      .sys_rst_n       (sys_rst_n),
      .hsi_clk         (hsi_clk),
      .csi_clk         (csi_clk),
      .hse_clk         (hse_clk),
      .pll1_p_clk      (pll1_p_clk),
      .sys_clk_sw      (sys_clk_sw),
      .d1cpre          (d1cpre),
      .d1ppre          (d1ppre),
      .hpre            (hpre),
      .d2ppre1         (d2ppre1),
      .d2ppre2         (d2ppre2),
      .d3ppre          (d3ppre),
      .timpre          (timpre),
      .hrtimsel        (hrtimsel),
      .c2_sleep        (c2_sleep),
      .c2_deepsleep    (c2_deepsleep),
      .c1_sleep        (c1_sleep),
      .c1_deepsleep    (c1_deepsleep),
      .d1_clk_arcg_en  (d1_clk_arcg_en),
      .d2_clk_arcg_en  (d2_clk_arcg_en),
      .cpu1_clk_arcg_en(cpu1_clk_arcg_en),
      .cpu2_clk_arcg_en(cpu2_clk_arcg_en),
      .sys_clk_arcg_en (sys_clk_arcg_en),
      .rcc_d1_stop     (rcc_d1_stop),
      .rcc_d2_stop     (rcc_d2_stop),
      .rcc_sys_stop    (rcc_sys_stop),

      .rcc_c2_clk               (rcc_c2_clk),
      .rcc_fclk_c2              (rcc_fclk_c2),
      .rcc_c2_systick_clk       (rcc_c2_systick_clk),
      .rcc_c1_clk               (rcc_c1_clk),
      .rcc_fclk_c1              (rcc_fclk_c1),
      .rcc_c1_systick_clk       (rcc_c1_systick_clk),
      .rcc_axibridge_d1_clk     (rcc_axibridge_d1_clk),
      .rcc_ahb3bridge_d1_clk    (rcc_ahb3bridge_d1_clk),
      .rcc_apb3bridge_d1_clk    (rcc_apb3bridge_d1_clk),
      .rcc_ahb1bridge_d2_clk    (rcc_ahb1bridge_d2_clk),
      .rcc_ahb2bridge_d2_clk    (rcc_ahb2bridge_d2_clk),
      .rcc_apb1bridge_d2_clk    (rcc_apb1bridge_d2_clk),
      .rcc_apb2bridge_d2_clk    (rcc_apb2bridge_d2_clk),
      .rcc_ahb4bridge_d3_clk    (rcc_ahb4bridge_d3_clk),
      .rcc_apb4bridge_d3_clk    (rcc_apb4bridge_d3_clk),
      .rcc_timx_ker_clk         (rcc_timx_ker_clk),
      .rcc_timy_ker_clk         (rcc_timy_ker_clk),
      .rcc_hrtimer_prescalar_clk(rcc_hrtimer_prescalar_clk),
      .sys_d1cpre_clk           (sys_d1cpre_clk),
      .sys_hpre_clk             (sys_hpre_clk),
      .sys_clk                  (sys_clk),
      .sys_clk_pre              (sys_clk_pre)
  );
  rcc_eth_ker_clk_ctrl u_rcc_eth_ker_clk_ctrl (
      .pad_rcc_eth_mii_tx_clk(pad_rcc_eth_mii_tx_clk),
      .pad_rcc_eth_mii_rx_clk(pad_rcc_eth_mii_rx_clk),
      .eth_rcc_fes           (eth_rcc_fes),
      .eth_rcc_epis_2        (eth_rcc_epis_2),
      .rst_n                 (sys_rst_n),
      .c1_sleep              (c1_sleep),
      .c1_deepsleep          (c1_deepsleep),
      .c2_sleep              (c2_sleep),
      .c2_deepsleep          (c2_deepsleep),
      .rcc_c1_eth1rx_en      (rcc_c1_eth1rx_en),
      .rcc_c2_eth1rx_en      (rcc_c2_eth1rx_en),
      .rcc_c1_eth1rx_lpen    (rcc_c1_eth1rx_lpen),
      .rcc_c2_eth1rx_lpen    (rcc_c2_eth1rx_lpen),
      .rcc_c1_eth1tx_en      (rcc_c1_eth1tx_en),
      .rcc_c2_eth1tx_en      (rcc_c2_eth1tx_en),
      .rcc_c1_eth1tx_lpen    (rcc_c1_eth1tx_lpen),
      .rcc_c2_eth1tx_lpen    (rcc_c2_eth1tx_lpen),

      .rcc_eth_mii_tx_clk  (rcc_eth_mii_tx_clk),
      .rcc_eth_mii_rx_clk  (rcc_eth_mii_rx_clk),
      .rcc_eth_rmii_ref_clk(rcc_eth_rmii_ref_clk)
  );

  rcc_per_clk_control u_rcc_per_clk_control (
      .sys_rst_n               (sys_rst_n),
      .rcc_axibridge_d1_clk    (rcc_axibridge_d1_clk),
      .rcc_ahb3bridge_d1_clk   (rcc_ahb3bridge_d1_clk),
      .rcc_apb3bridge_d1_clk   (rcc_apb3bridge_d1_clk),
      .rcc_ahb1bridge_d2_clk   (rcc_ahb1bridge_d2_clk),
      .rcc_ahb2bridge_d2_clk   (rcc_ahb2bridge_d2_clk),
      .rcc_apb1bridge_d2_clk   (rcc_apb1bridge_d2_clk),
      .rcc_apb2bridge_d2_clk   (rcc_apb2bridge_d2_clk),
      .rcc_ahb4bridge_d3_clk   (rcc_ahb4bridge_d3_clk),
      .rcc_apb4bridge_d3_clk   (rcc_apb4bridge_d3_clk),
      .pll1_q_clk              (pll1_q_clk),
      .pll2_p_clk              (pll2_p_clk),
      .pll2_q_clk              (pll2_q_clk),
      .pll2_r_clk              (pll2_r_clk),
      .pll3_p_clk              (pll3_p_clk),
      .pll3_q_clk              (pll3_q_clk),
      .pll3_r_clk              (pll3_r_clk),
      .sys_clk                 (sys_clk),
      .hse_clk                 (hse_clk),
      .hsi_ker_clk             (hsi_ker_clk),
      .csi_ker_clk             (csi_ker_clk),
      .hsi48_clk               (hsi48_clk),
      .lse_clk                 (lse_clk),
      .lsi_clk                 (lsi_clk),
      .per_clk                 (per_clk),
      .I2S_clk_IN              (I2S_clk_IN),
      .USB_PHY1                (USB_PHY1),
      .c1_sleep                (c1_sleep),
      .c1_deepsleep            (c1_deepsleep),
      .c2_sleep                (c2_sleep),
      .c2_deepsleep            (c2_deepsleep),
      .d3_deepsleep            (d3_deepsleep),
      .rcc_flash_arcg_clk_en   (rcc_flash_arcg_clk_en),
      .rcc_c2_flash_en         (rcc_c2_flash_en),
      .rcc_c1_flash_lpen       (rcc_c1_flash_lpen),
      .rcc_c2_flash_lpen       (rcc_c2_flash_lpen),
      .rcc_qspi_arcg_clk_en    (rcc_qspi_arcg_clk_en),
      .rcc_c1_qspi_en          (rcc_c1_qspi_en),
      .rcc_c2_qspi_en          (rcc_c2_qspi_en),
      .rcc_c1_qspi_lpen        (rcc_c1_qspi_lpen),
      .rcc_c2_qspi_lpen        (rcc_c2_qspi_lpen),
      .rcc_axisram_arcg_clk_en (rcc_axisram_arcg_clk_en),
      .rcc_c2_axisram_en       (rcc_c2_axisram_en),
      .rcc_c1_axisram_lpen     (rcc_c1_axisram_lpen),
      .rcc_c2_axisram_lpen     (rcc_c2_axisram_lpen),
      .rcc_fmc_arcg_clk_en     (rcc_fmc_arcg_clk_en),
      .rcc_c1_fmc_en           (rcc_c1_fmc_en),
      .rcc_c2_fmc_en           (rcc_c2_fmc_en),
      .rcc_c1_fmc_lpen         (rcc_c1_fmc_lpen),
      .rcc_c2_fmc_lpen         (rcc_c2_fmc_lpen),
      .rcc_dma2d_arcg_clk_en   (rcc_dma2d_arcg_clk_en),
      .rcc_c1_dma2d_en         (rcc_c1_dma2d_en),
      .rcc_c2_dma2d_en         (rcc_c2_dma2d_en),
      .rcc_c1_dma2d_lpen       (rcc_c1_dma2d_lpen),
      .rcc_c2_dma2d_lpen       (rcc_c2_dma2d_lpen),
      .rcc_mdma_arcg_clk_en    (rcc_mdma_arcg_clk_en),
      .rcc_c1_mdma_en          (rcc_c1_mdma_en),
      .rcc_c2_mdma_en          (rcc_c2_mdma_en),
      .rcc_c1_mdma_lpen        (rcc_c1_mdma_lpen),
      .rcc_c2_mdma_lpen        (rcc_c2_mdma_lpen),
      .rcc_ltdc_arcg_clk_en    (rcc_ltdc_arcg_clk_en),
      .rcc_c1_ltdc_en          (rcc_c1_ltdc_en),
      .rcc_c2_ltdc_en          (rcc_c2_ltdc_en),
      .rcc_c1_ltdc_lpen        (rcc_c1_ltdc_lpen),
      .rcc_c2_ltdc_lpen        (rcc_c2_ltdc_lpen),
      .rcc_ramecc1_arcg_clk_en (rcc_ramecc1_arcg_clk_en),
      .rcc_gpv_arcg_clk_en     (rcc_gpv_arcg_clk_en),
      .rcc_itcm_arcg_clk_en    (rcc_itcm_arcg_clk_en),
      .rcc_c2_itcm_en          (rcc_c2_itcm_en),
      .rcc_c1_itcm_lpen        (rcc_c1_itcm_lpen),
      .rcc_c2_itcm_lpen        (rcc_c2_itcm_lpen),
      .rcc_dtcm2_arcg_clk_en   (rcc_dtcm2_arcg_clk_en),
      .rcc_c2_dtcm2_en         (rcc_c2_dtcm2_en),
      .rcc_c1_dtcm2_lpen       (rcc_c1_dtcm2_lpen),
      .rcc_c2_dtcm2_lpen       (rcc_c2_dtcm2_lpen),
      .rcc_dtcm1_arcg_clk_en   (rcc_dtcm1_arcg_clk_en),
      .rcc_c2_dtcm1_en         (rcc_c2_dtcm1_en),
      .rcc_c1_dtcm1_lpen       (rcc_c1_dtcm1_lpen),
      .rcc_c2_dtcm1_lpen       (rcc_c2_dtcm1_lpen),
      .rcc_jpgdec_arcg_clk_en  (rcc_jpgdec_arcg_clk_en),
      .rcc_c1_jpgdec_en        (rcc_c1_jpgdec_en),
      .rcc_c2_jpgdec_en        (rcc_c2_jpgdec_en),
      .rcc_c1_jpgdec_lpen      (rcc_c1_jpgdec_lpen),
      .rcc_c2_jpgdec_lpen      (rcc_c2_jpgdec_lpen),
      .rcc_sdmmc1_arcg_clk_en  (rcc_sdmmc1_arcg_clk_en),
      .rcc_c1_sdmmc1_en        (rcc_c1_sdmmc1_en),
      .rcc_c2_sdmmc1_en        (rcc_c2_sdmmc1_en),
      .rcc_c1_sdmmc1_lpen      (rcc_c1_sdmmc1_lpen),
      .rcc_c2_sdmmc1_lpen      (rcc_c2_sdmmc1_lpen),
      .rcc_wwdg1_arcg_clk_en   (rcc_wwdg1_arcg_clk_en),
      .rcc_c1_wwdg1_en         (rcc_c1_wwdg1_en),
      .rcc_c2_wwdg1_en         (rcc_c2_wwdg1_en),
      .rcc_c1_wwdg1_lpen       (rcc_c1_wwdg1_lpen),
      .rcc_c2_wwdg1_lpen       (rcc_c2_wwdg1_lpen),
      .rcc_usb2ulpi_arcg_clk_en(rcc_usb2ulpi_arcg_clk_en),
      .rcc_c1_usb2ulpi_en      (rcc_c1_usb2ulpi_en),
      .rcc_c2_usb2ulpi_en      (rcc_c2_usb2ulpi_en),
      .rcc_c1_usb2ulpi_lpen    (rcc_c1_usb2ulpi_lpen),
      .rcc_c2_usb2ulpi_lpen    (rcc_c2_usb2ulpi_lpen),
      .rcc_usb2otg_arcg_clk_en (rcc_usb2otg_arcg_clk_en),
      .rcc_c1_usb2otg_en       (rcc_c1_usb2otg_en),
      .rcc_c2_usb2otg_en       (rcc_c2_usb2otg_en),
      .rcc_c1_usb2otg_lpen     (rcc_c1_usb2otg_lpen),
      .rcc_c2_usb2otg_lpen     (rcc_c2_usb2otg_lpen),
      .rcc_usb1ulpi_arcg_clk_en(rcc_usb1ulpi_arcg_clk_en),
      .rcc_c1_usb1ulpi_en      (rcc_c1_usb1ulpi_en),
      .rcc_c2_usb1ulpi_en      (rcc_c2_usb1ulpi_en),
      .rcc_c1_usb1ulpi_lpen    (rcc_c1_usb1ulpi_lpen),
      .rcc_c2_usb1ulpi_lpen    (rcc_c2_usb1ulpi_lpen),
      .rcc_usb1otg_arcg_clk_en (rcc_usb1otg_arcg_clk_en),
      .rcc_c1_usb1otg_en       (rcc_c1_usb1otg_en),
      .rcc_c2_usb1otg_en       (rcc_c2_usb1otg_en),
      .rcc_c1_usb1otg_lpen     (rcc_c1_usb1otg_lpen),
      .rcc_c2_usb1otg_lpen     (rcc_c2_usb1otg_lpen),
      .rcc_eth1rx_arcg_clk_en  (rcc_eth1rx_arcg_clk_en),
      .rcc_c1_eth1rx_en        (rcc_c1_eth1rx_en),
      .rcc_c2_eth1rx_en        (rcc_c2_eth1rx_en),
      .rcc_c1_eth1rx_lpen      (rcc_c1_eth1rx_lpen),
      .rcc_c2_eth1rx_lpen      (rcc_c2_eth1rx_lpen),
      .rcc_eth1tx_arcg_clk_en  (rcc_eth1tx_arcg_clk_en),
      .rcc_c1_eth1tx_en        (rcc_c1_eth1tx_en),
      .rcc_c2_eth1tx_en        (rcc_c2_eth1tx_en),
      .rcc_c1_eth1tx_lpen      (rcc_c1_eth1tx_lpen),
      .rcc_c2_eth1tx_lpen      (rcc_c2_eth1tx_lpen),
      .rcc_eth1mac_arcg_clk_en (rcc_eth1mac_arcg_clk_en),
      .rcc_c1_eth1mac_en       (rcc_c1_eth1mac_en),
      .rcc_c2_eth1mac_en       (rcc_c2_eth1mac_en),
      .rcc_c1_eth1mac_lpen     (rcc_c1_eth1mac_lpen),
      .rcc_c2_eth1mac_lpen     (rcc_c2_eth1mac_lpen),
      .rcc_adc12_arcg_clk_en   (rcc_adc12_arcg_clk_en),
      .rcc_c1_adc12_en         (rcc_c1_adc12_en),
      .rcc_c2_adc12_en         (rcc_c2_adc12_en),
      .rcc_c1_adc12_lpen       (rcc_c1_adc12_lpen),
      .rcc_c2_adc12_lpen       (rcc_c2_adc12_lpen),
      .rcc_dma2_arcg_clk_en    (rcc_dma2_arcg_clk_en),
      .rcc_c1_dma2_en          (rcc_c1_dma2_en),
      .rcc_c2_dma2_en          (rcc_c2_dma2_en),
      .rcc_c1_dma2_lpen        (rcc_c1_dma2_lpen),
      .rcc_c2_dma2_lpen        (rcc_c2_dma2_lpen),
      .rcc_dma1_arcg_clk_en    (rcc_dma1_arcg_clk_en),
      .rcc_c1_dma1_en          (rcc_c1_dma1_en),
      .rcc_c2_dma1_en          (rcc_c2_dma1_en),
      .rcc_c1_dma1_lpen        (rcc_c1_dma1_lpen),
      .rcc_c2_dma1_lpen        (rcc_c2_dma1_lpen),
      .rcc_sram3_arcg_clk_en   (rcc_sram3_arcg_clk_en),
      .rcc_c1_sram3_en         (rcc_c1_sram3_en),
      .rcc_c1_sram3_lpen       (rcc_c1_sram3_lpen),
      .rcc_c2_sram3_lpen       (rcc_c2_sram3_lpen),
      .rcc_sram2_arcg_clk_en   (rcc_sram2_arcg_clk_en),
      .rcc_c1_sram2_en         (rcc_c1_sram2_en),
      .rcc_c1_sram2_lpen       (rcc_c1_sram2_lpen),
      .rcc_c2_sram2_lpen       (rcc_c2_sram2_lpen),
      .rcc_sram1_arcg_clk_en   (rcc_sram1_arcg_clk_en),
      .rcc_c1_sram1_en         (rcc_c1_sram1_en),
      .rcc_c1_sram1_lpen       (rcc_c1_sram1_lpen),
      .rcc_c2_sram1_lpen       (rcc_c2_sram1_lpen),
      .rcc_sdmmc2_arcg_clk_en  (rcc_sdmmc2_arcg_clk_en),
      .rcc_c1_sdmmc2_en        (rcc_c1_sdmmc2_en),
      .rcc_c2_sdmmc2_en        (rcc_c2_sdmmc2_en),
      .rcc_c1_sdmmc2_lpen      (rcc_c1_sdmmc2_lpen),
      .rcc_c2_sdmmc2_lpen      (rcc_c2_sdmmc2_lpen),
      .rcc_rng_arcg_clk_en     (rcc_rng_arcg_clk_en),
      .rcc_c1_rng_en           (rcc_c1_rng_en),
      .rcc_c2_rng_en           (rcc_c2_rng_en),
      .rcc_c1_rng_lpen         (rcc_c1_rng_lpen),
      .rcc_c2_rng_lpen         (rcc_c2_rng_lpen),
      .rcc_hash_arcg_clk_en    (rcc_hash_arcg_clk_en),
      .rcc_c1_hash_en          (rcc_c1_hash_en),
      .rcc_c2_hash_en          (rcc_c2_hash_en),
      .rcc_c1_hash_lpen        (rcc_c1_hash_lpen),
      .rcc_c2_hash_lpen        (rcc_c2_hash_lpen),
      .rcc_crypt_arcg_clk_en   (rcc_crypt_arcg_clk_en),
      .rcc_c1_crypt_en         (rcc_c1_crypt_en),
      .rcc_c2_crypt_en         (rcc_c2_crypt_en),
      .rcc_c1_crypt_lpen       (rcc_c1_crypt_lpen),
      .rcc_c2_crypt_lpen       (rcc_c2_crypt_lpen),
      .rcc_dcmi_arcg_clk_en    (rcc_dcmi_arcg_clk_en),
      .rcc_c1_dcmi_en          (rcc_c1_dcmi_en),
      .rcc_c2_dcmi_en          (rcc_c2_dcmi_en),
      .rcc_c1_dcmi_lpen        (rcc_c1_dcmi_lpen),
      .rcc_c2_dcmi_lpen        (rcc_c2_dcmi_lpen),
      .rcc_ramecc2_arcg_clk_en (rcc_ramecc2_arcg_clk_en),
      .rcc_uart8_arcg_clk_en   (rcc_uart8_arcg_clk_en),
      .rcc_c1_uart8_en         (rcc_c1_uart8_en),
      .rcc_c2_uart8_en         (rcc_c2_uart8_en),
      .rcc_c1_uart8_lpen       (rcc_c1_uart8_lpen),
      .rcc_c2_uart8_lpen       (rcc_c2_uart8_lpen),
      .uart8_ker_clk_req       (uart8_ker_clk_req),
      .rcc_uart7_arcg_clk_en   (rcc_uart7_arcg_clk_en),
      .rcc_c1_uart7_en         (rcc_c1_uart7_en),
      .rcc_c2_uart7_en         (rcc_c2_uart7_en),
      .rcc_c1_uart7_lpen       (rcc_c1_uart7_lpen),
      .rcc_c2_uart7_lpen       (rcc_c2_uart7_lpen),
      .uart7_ker_clk_req       (uart7_ker_clk_req),
      .rcc_dac12_arcg_clk_en   (rcc_dac12_arcg_clk_en),
      .rcc_c1_dac12_en         (rcc_c1_dac12_en),
      .rcc_c2_dac12_en         (rcc_c2_dac12_en),
      .rcc_c1_dac12_lpen       (rcc_c1_dac12_lpen),
      .rcc_c2_dac12_lpen       (rcc_c2_dac12_lpen),
      .rcc_hdmicec_arcg_clk_en (rcc_hdmicec_arcg_clk_en),
      .rcc_c1_hdmicec_en       (rcc_c1_hdmicec_en),
      .rcc_c2_hdmicec_en       (rcc_c2_hdmicec_en),
      .rcc_c1_hdmicec_lpen     (rcc_c1_hdmicec_lpen),
      .rcc_c2_hdmicec_lpen     (rcc_c2_hdmicec_lpen),
      .rcc_i2c3_arcg_clk_en    (rcc_i2c3_arcg_clk_en),
      .rcc_c1_i2c3_en          (rcc_c1_i2c3_en),
      .rcc_c2_i2c3_en          (rcc_c2_i2c3_en),
      .rcc_c1_i2c3_lpen        (rcc_c1_i2c3_lpen),
      .rcc_c2_i2c3_lpen        (rcc_c2_i2c3_lpen),
      .i2c3_ker_clk_req        (i2c3_ker_clk_req),
      .rcc_i2c2_arcg_clk_en    (rcc_i2c2_arcg_clk_en),
      .rcc_c1_i2c2_en          (rcc_c1_i2c2_en),
      .rcc_c2_i2c2_en          (rcc_c2_i2c2_en),
      .rcc_c1_i2c2_lpen        (rcc_c1_i2c2_lpen),
      .rcc_c2_i2c2_lpen        (rcc_c2_i2c2_lpen),
      .i2c2_ker_clk_req        (i2c2_ker_clk_req),
      .rcc_i2c1_arcg_clk_en    (rcc_i2c1_arcg_clk_en),
      .rcc_c1_i2c1_en          (rcc_c1_i2c1_en),
      .rcc_c2_i2c1_en          (rcc_c2_i2c1_en),
      .rcc_c1_i2c1_lpen        (rcc_c1_i2c1_lpen),
      .rcc_c2_i2c1_lpen        (rcc_c2_i2c1_lpen),
      .i2c1_ker_clk_req        (i2c1_ker_clk_req),
      .rcc_uart5_arcg_clk_en   (rcc_uart5_arcg_clk_en),
      .rcc_c1_uart5_en         (rcc_c1_uart5_en),
      .rcc_c2_uart5_en         (rcc_c2_uart5_en),
      .rcc_c1_uart5_lpen       (rcc_c1_uart5_lpen),
      .rcc_c2_uart5_lpen       (rcc_c2_uart5_lpen),
      .uart5_ker_clk_req       (uart5_ker_clk_req),
      .rcc_uart4_arcg_clk_en   (rcc_uart4_arcg_clk_en),
      .rcc_c1_uart4_en         (rcc_c1_uart4_en),
      .rcc_c2_uart4_en         (rcc_c2_uart4_en),
      .rcc_c1_uart4_lpen       (rcc_c1_uart4_lpen),
      .rcc_c2_uart4_lpen       (rcc_c2_uart4_lpen),
      .uart4_ker_clk_req       (uart4_ker_clk_req),
      .rcc_usart3_arcg_clk_en  (rcc_usart3_arcg_clk_en),
      .rcc_c1_usart3_en        (rcc_c1_usart3_en),
      .rcc_c2_usart3_en        (rcc_c2_usart3_en),
      .rcc_c1_usart3_lpen      (rcc_c1_usart3_lpen),
      .rcc_c2_usart3_lpen      (rcc_c2_usart3_lpen),
      .usart3_ker_clk_req      (usart3_ker_clk_req),
      .rcc_usart2_arcg_clk_en  (rcc_usart2_arcg_clk_en),
      .rcc_c1_usart2_en        (rcc_c1_usart2_en),
      .rcc_c2_usart2_en        (rcc_c2_usart2_en),
      .rcc_c1_usart2_lpen      (rcc_c1_usart2_lpen),
      .rcc_c2_usart2_lpen      (rcc_c2_usart2_lpen),
      .usart2_ker_clk_req      (usart2_ker_clk_req),
      .rcc_spdifrx_arcg_clk_en (rcc_spdifrx_arcg_clk_en),
      .rcc_c1_spdifrx_en       (rcc_c1_spdifrx_en),
      .rcc_c2_spdifrx_en       (rcc_c2_spdifrx_en),
      .rcc_c1_spdifrx_lpen     (rcc_c1_spdifrx_lpen),
      .rcc_c2_spdifrx_lpen     (rcc_c2_spdifrx_lpen),
      .rcc_spi3_arcg_clk_en    (rcc_spi3_arcg_clk_en),
      .rcc_c1_spi3_en          (rcc_c1_spi3_en),
      .rcc_c2_spi3_en          (rcc_c2_spi3_en),
      .rcc_c1_spi3_lpen        (rcc_c1_spi3_lpen),
      .rcc_c2_spi3_lpen        (rcc_c2_spi3_lpen),
      .rcc_spi2_arcg_clk_en    (rcc_spi2_arcg_clk_en),
      .rcc_c1_spi2_en          (rcc_c1_spi2_en),
      .rcc_c2_spi2_en          (rcc_c2_spi2_en),
      .rcc_c1_spi2_lpen        (rcc_c1_spi2_lpen),
      .rcc_c2_spi2_lpen        (rcc_c2_spi2_lpen),
      .rcc_wwdg2_arcg_clk_en   (rcc_wwdg2_arcg_clk_en),
      .rcc_c1_wwdg2_en         (rcc_c1_wwdg2_en),
      .rcc_c2_wwdg2_en         (rcc_c2_wwdg2_en),
      .rcc_c1_wwdg2_lpen       (rcc_c1_wwdg2_lpen),
      .rcc_c2_wwdg2_lpen       (rcc_c2_wwdg2_lpen),
      .rcc_lptim1_arcg_clk_en  (rcc_lptim1_arcg_clk_en),
      .rcc_c1_lptim1_en        (rcc_c1_lptim1_en),
      .rcc_c2_lptim1_en        (rcc_c2_lptim1_en),
      .rcc_c1_lptim1_lpen      (rcc_c1_lptim1_lpen),
      .rcc_c2_lptim1_lpen      (rcc_c2_lptim1_lpen),
      .rcc_tim14_arcg_clk_en   (rcc_tim14_arcg_clk_en),
      .rcc_c1_tim14_en         (rcc_c1_tim14_en),
      .rcc_c2_tim14_en         (rcc_c2_tim14_en),
      .rcc_c1_tim14_lpen       (rcc_c1_tim14_lpen),
      .rcc_c2_tim14_lpen       (rcc_c2_tim14_lpen),
      .rcc_tim13_arcg_clk_en   (rcc_tim13_arcg_clk_en),
      .rcc_c1_tim13_en         (rcc_c1_tim13_en),
      .rcc_c2_tim13_en         (rcc_c2_tim13_en),
      .rcc_c1_tim13_lpen       (rcc_c1_tim13_lpen),
      .rcc_c2_tim13_lpen       (rcc_c2_tim13_lpen),
      .rcc_tim12_arcg_clk_en   (rcc_tim12_arcg_clk_en),
      .rcc_c1_tim12_en         (rcc_c1_tim12_en),
      .rcc_c2_tim12_en         (rcc_c2_tim12_en),
      .rcc_c1_tim12_lpen       (rcc_c1_tim12_lpen),
      .rcc_c2_tim12_lpen       (rcc_c2_tim12_lpen),
      .rcc_tim7_arcg_clk_en    (rcc_tim7_arcg_clk_en),
      .rcc_c1_tim7_en          (rcc_c1_tim7_en),
      .rcc_c2_tim7_en          (rcc_c2_tim7_en),
      .rcc_c1_tim7_lpen        (rcc_c1_tim7_lpen),
      .rcc_c2_tim7_lpen        (rcc_c2_tim7_lpen),
      .rcc_tim6_arcg_clk_en    (rcc_tim6_arcg_clk_en),
      .rcc_c1_tim6_en          (rcc_c1_tim6_en),
      .rcc_c2_tim6_en          (rcc_c2_tim6_en),
      .rcc_c1_tim6_lpen        (rcc_c1_tim6_lpen),
      .rcc_c2_tim6_lpen        (rcc_c2_tim6_lpen),
      .rcc_tim5_arcg_clk_en    (rcc_tim5_arcg_clk_en),
      .rcc_c1_tim5_en          (rcc_c1_tim5_en),
      .rcc_c2_tim5_en          (rcc_c2_tim5_en),
      .rcc_c1_tim5_lpen        (rcc_c1_tim5_lpen),
      .rcc_c2_tim5_lpen        (rcc_c2_tim5_lpen),
      .rcc_tim4_arcg_clk_en    (rcc_tim4_arcg_clk_en),
      .rcc_c1_tim4_en          (rcc_c1_tim4_en),
      .rcc_c2_tim4_en          (rcc_c2_tim4_en),
      .rcc_c1_tim4_lpen        (rcc_c1_tim4_lpen),
      .rcc_c2_tim4_lpen        (rcc_c2_tim4_lpen),
      .rcc_tim3_arcg_clk_en    (rcc_tim3_arcg_clk_en),
      .rcc_c1_tim3_en          (rcc_c1_tim3_en),
      .rcc_c2_tim3_en          (rcc_c2_tim3_en),
      .rcc_c1_tim3_lpen        (rcc_c1_tim3_lpen),
      .rcc_c2_tim3_lpen        (rcc_c2_tim3_lpen),
      .rcc_tim2_arcg_clk_en    (rcc_tim2_arcg_clk_en),
      .rcc_c1_tim2_en          (rcc_c1_tim2_en),
      .rcc_c2_tim2_en          (rcc_c2_tim2_en),
      .rcc_c1_tim2_lpen        (rcc_c1_tim2_lpen),
      .rcc_c2_tim2_lpen        (rcc_c2_tim2_lpen),
      .rcc_fdcan_arcg_clk_en   (rcc_fdcan_arcg_clk_en),
      .rcc_c1_fdcan_en         (rcc_c1_fdcan_en),
      .rcc_c2_fdcan_en         (rcc_c2_fdcan_en),
      .rcc_c1_fdcan_lpen       (rcc_c1_fdcan_lpen),
      .rcc_c2_fdcan_lpen       (rcc_c2_fdcan_lpen),
      .rcc_mdios_arcg_clk_en   (rcc_mdios_arcg_clk_en),
      .rcc_c1_mdios_en         (rcc_c1_mdios_en),
      .rcc_c2_mdios_en         (rcc_c2_mdios_en),
      .rcc_c1_mdios_lpen       (rcc_c1_mdios_lpen),
      .rcc_c2_mdios_lpen       (rcc_c2_mdios_lpen),
      .rcc_opamp_arcg_clk_en   (rcc_opamp_arcg_clk_en),
      .rcc_c1_opamp_en         (rcc_c1_opamp_en),
      .rcc_c2_opamp_en         (rcc_c2_opamp_en),
      .rcc_c1_opamp_lpen       (rcc_c1_opamp_lpen),
      .rcc_c2_opamp_lpen       (rcc_c2_opamp_lpen),
      .rcc_swpmi_arcg_clk_en   (rcc_swpmi_arcg_clk_en),
      .rcc_c1_swpmi_en         (rcc_c1_swpmi_en),
      .rcc_c2_swpmi_en         (rcc_c2_swpmi_en),
      .rcc_c1_swpmi_lpen       (rcc_c1_swpmi_lpen),
      .rcc_c2_swpmi_lpen       (rcc_c2_swpmi_lpen),
      .rcc_crs_arcg_clk_en     (rcc_crs_arcg_clk_en),
      .rcc_c1_crs_en           (rcc_c1_crs_en),
      .rcc_c2_crs_en           (rcc_c2_crs_en),
      .rcc_c1_crs_lpen         (rcc_c1_crs_lpen),
      .rcc_c2_crs_lpen         (rcc_c2_crs_lpen),
      .rcc_hrtim_arcg_clk_en   (rcc_hrtim_arcg_clk_en),
      .rcc_c1_hrtim_en         (rcc_c1_hrtim_en),
      .rcc_c2_hrtim_en         (rcc_c2_hrtim_en),
      .rcc_c1_hrtim_lpen       (rcc_c1_hrtim_lpen),
      .rcc_c2_hrtim_lpen       (rcc_c2_hrtim_lpen),
      .rcc_dfsdm1_arcg_clk_en  (rcc_dfsdm1_arcg_clk_en),
      .rcc_c1_dfsdm1_en        (rcc_c1_dfsdm1_en),
      .rcc_c2_dfsdm1_en        (rcc_c2_dfsdm1_en),
      .rcc_c1_dfsdm1_lpen      (rcc_c1_dfsdm1_lpen),
      .rcc_c2_dfsdm1_lpen      (rcc_c2_dfsdm1_lpen),
      .rcc_sai3_arcg_clk_en    (rcc_sai3_arcg_clk_en),
      .rcc_c1_sai3_en          (rcc_c1_sai3_en),
      .rcc_c2_sai3_en          (rcc_c2_sai3_en),
      .rcc_c1_sai3_lpen        (rcc_c1_sai3_lpen),
      .rcc_c2_sai3_lpen        (rcc_c2_sai3_lpen),
      .rcc_sai2_arcg_clk_en    (rcc_sai2_arcg_clk_en),
      .rcc_c1_sai2_en          (rcc_c1_sai2_en),
      .rcc_c2_sai2_en          (rcc_c2_sai2_en),
      .rcc_c1_sai2_lpen        (rcc_c1_sai2_lpen),
      .rcc_c2_sai2_lpen        (rcc_c2_sai2_lpen),
      .rcc_sai1_arcg_clk_en    (rcc_sai1_arcg_clk_en),
      .rcc_c1_sai1_en          (rcc_c1_sai1_en),
      .rcc_c2_sai1_en          (rcc_c2_sai1_en),
      .rcc_c1_sai1_lpen        (rcc_c1_sai1_lpen),
      .rcc_c2_sai1_lpen        (rcc_c2_sai1_lpen),
      .rcc_spi5_arcg_clk_en    (rcc_spi5_arcg_clk_en),
      .rcc_c1_spi5_en          (rcc_c1_spi5_en),
      .rcc_c2_spi5_en          (rcc_c2_spi5_en),
      .rcc_c1_spi5_lpen        (rcc_c1_spi5_lpen),
      .rcc_c2_spi5_lpen        (rcc_c2_spi5_lpen),
      .rcc_tim17_arcg_clk_en   (rcc_tim17_arcg_clk_en),
      .rcc_c1_tim17_en         (rcc_c1_tim17_en),
      .rcc_c2_tim17_en         (rcc_c2_tim17_en),
      .rcc_c1_tim17_lpen       (rcc_c1_tim17_lpen),
      .rcc_c2_tim17_lpen       (rcc_c2_tim17_lpen),
      .rcc_tim16_arcg_clk_en   (rcc_tim16_arcg_clk_en),
      .rcc_c1_tim16_en         (rcc_c1_tim16_en),
      .rcc_c2_tim16_en         (rcc_c2_tim16_en),
      .rcc_c1_tim16_lpen       (rcc_c1_tim16_lpen),
      .rcc_c2_tim16_lpen       (rcc_c2_tim16_lpen),
      .rcc_tim15_arcg_clk_en   (rcc_tim15_arcg_clk_en),
      .rcc_c1_tim15_en         (rcc_c1_tim15_en),
      .rcc_c2_tim15_en         (rcc_c2_tim15_en),
      .rcc_c1_tim15_lpen       (rcc_c1_tim15_lpen),
      .rcc_c2_tim15_lpen       (rcc_c2_tim15_lpen),
      .rcc_spi4_arcg_clk_en    (rcc_spi4_arcg_clk_en),
      .rcc_c1_spi4_en          (rcc_c1_spi4_en),
      .rcc_c2_spi4_en          (rcc_c2_spi4_en),
      .rcc_c1_spi4_lpen        (rcc_c1_spi4_lpen),
      .rcc_c2_spi4_lpen        (rcc_c2_spi4_lpen),
      .rcc_spi1_arcg_clk_en    (rcc_spi1_arcg_clk_en),
      .rcc_c1_spi1_en          (rcc_c1_spi1_en),
      .rcc_c2_spi1_en          (rcc_c2_spi1_en),
      .rcc_c1_spi1_lpen        (rcc_c1_spi1_lpen),
      .rcc_c2_spi1_lpen        (rcc_c2_spi1_lpen),
      .rcc_usart6_arcg_clk_en  (rcc_usart6_arcg_clk_en),
      .rcc_c1_usart6_en        (rcc_c1_usart6_en),
      .rcc_c2_usart6_en        (rcc_c2_usart6_en),
      .rcc_c1_usart6_lpen      (rcc_c1_usart6_lpen),
      .rcc_c2_usart6_lpen      (rcc_c2_usart6_lpen),
      .usart6_ker_clk_req      (usart6_ker_clk_req),
      .rcc_usart1_arcg_clk_en  (rcc_usart1_arcg_clk_en),
      .rcc_c1_usart1_en        (rcc_c1_usart1_en),
      .rcc_c2_usart1_en        (rcc_c2_usart1_en),
      .rcc_c1_usart1_lpen      (rcc_c1_usart1_lpen),
      .rcc_c2_usart1_lpen      (rcc_c2_usart1_lpen),
      .usart1_ker_clk_req      (usart1_ker_clk_req),
      .rcc_tim8_arcg_clk_en    (rcc_tim8_arcg_clk_en),
      .rcc_c1_tim8_en          (rcc_c1_tim8_en),
      .rcc_c2_tim8_en          (rcc_c2_tim8_en),
      .rcc_c1_tim8_lpen        (rcc_c1_tim8_lpen),
      .rcc_c2_tim8_lpen        (rcc_c2_tim8_lpen),
      .rcc_tim1_arcg_clk_en    (rcc_tim1_arcg_clk_en),
      .rcc_c1_tim1_en          (rcc_c1_tim1_en),
      .rcc_c2_tim1_en          (rcc_c2_tim1_en),
      .rcc_c1_tim1_lpen        (rcc_c1_tim1_lpen),
      .rcc_c2_tim1_lpen        (rcc_c2_tim1_lpen),
      .rcc_sram4_arcg_clk_en   (rcc_sram4_arcg_clk_en),
      .rcc_c1_sram4_lpen       (rcc_c1_sram4_lpen),
      .rcc_c2_sram4_lpen       (rcc_c2_sram4_lpen),
      .rcc_sram4_amen          (rcc_sram4_amen),
      .rcc_bkpram_arcg_clk_en  (rcc_bkpram_arcg_clk_en),
      .rcc_c1_bkpram_en        (rcc_c1_bkpram_en),
      .rcc_c2_bkpram_en        (rcc_c2_bkpram_en),
      .rcc_c1_bkpram_lpen      (rcc_c1_bkpram_lpen),
      .rcc_c2_bkpram_lpen      (rcc_c2_bkpram_lpen),
      .rcc_bkpram_amen         (rcc_bkpram_amen),
      .rcc_ramecc3_arcg_clk_en (rcc_ramecc3_arcg_clk_en),
      .rcc_hsem_arcg_clk_en    (rcc_hsem_arcg_clk_en),
      .rcc_c1_hsem_en          (rcc_c1_hsem_en),
      .rcc_c2_hsem_en          (rcc_c2_hsem_en),
      .rcc_adc3_arcg_clk_en    (rcc_adc3_arcg_clk_en),
      .rcc_c1_adc3_en          (rcc_c1_adc3_en),
      .rcc_c2_adc3_en          (rcc_c2_adc3_en),
      .rcc_c1_adc3_lpen        (rcc_c1_adc3_lpen),
      .rcc_c2_adc3_lpen        (rcc_c2_adc3_lpen),
      .rcc_adc3_amen           (rcc_adc3_amen),
      .rcc_bdma_arcg_clk_en    (rcc_bdma_arcg_clk_en),
      .rcc_c1_bdma_en          (rcc_c1_bdma_en),
      .rcc_c2_bdma_en          (rcc_c2_bdma_en),
      .rcc_c1_bdma_lpen        (rcc_c1_bdma_lpen),
      .rcc_c2_bdma_lpen        (rcc_c2_bdma_lpen),
      .rcc_bdma_amen           (rcc_bdma_amen),
      .rcc_crc_arcg_clk_en     (rcc_crc_arcg_clk_en),
      .rcc_c1_crc_en           (rcc_c1_crc_en),
      .rcc_c2_crc_en           (rcc_c2_crc_en),
      .rcc_c1_crc_lpen         (rcc_c1_crc_lpen),
      .rcc_c2_crc_lpen         (rcc_c2_crc_lpen),
      .rcc_crc_amen            (rcc_crc_amen),
      .rcc_gpiok_arcg_clk_en   (rcc_gpiok_arcg_clk_en),
      .rcc_c1_gpiok_en         (rcc_c1_gpiok_en),
      .rcc_c2_gpiok_en         (rcc_c2_gpiok_en),
      .rcc_c1_gpiok_lpen       (rcc_c1_gpiok_lpen),
      .rcc_c2_gpiok_lpen       (rcc_c2_gpiok_lpen),
      .rcc_gpioj_arcg_clk_en   (rcc_gpioj_arcg_clk_en),
      .rcc_c1_gpioj_en         (rcc_c1_gpioj_en),
      .rcc_c2_gpioj_en         (rcc_c2_gpioj_en),
      .rcc_c1_gpioj_lpen       (rcc_c1_gpioj_lpen),
      .rcc_c2_gpioj_lpen       (rcc_c2_gpioj_lpen),
      .rcc_gpioi_arcg_clk_en   (rcc_gpioi_arcg_clk_en),
      .rcc_c1_gpioi_en         (rcc_c1_gpioi_en),
      .rcc_c2_gpioi_en         (rcc_c2_gpioi_en),
      .rcc_c1_gpioi_lpen       (rcc_c1_gpioi_lpen),
      .rcc_c2_gpioi_lpen       (rcc_c2_gpioi_lpen),
      .rcc_gpioh_arcg_clk_en   (rcc_gpioh_arcg_clk_en),
      .rcc_c1_gpioh_en         (rcc_c1_gpioh_en),
      .rcc_c2_gpioh_en         (rcc_c2_gpioh_en),
      .rcc_c1_gpioh_lpen       (rcc_c1_gpioh_lpen),
      .rcc_c2_gpioh_lpen       (rcc_c2_gpioh_lpen),
      .rcc_gpiog_arcg_clk_en   (rcc_gpiog_arcg_clk_en),
      .rcc_c1_gpiog_en         (rcc_c1_gpiog_en),
      .rcc_c2_gpiog_en         (rcc_c2_gpiog_en),
      .rcc_c1_gpiog_lpen       (rcc_c1_gpiog_lpen),
      .rcc_c2_gpiog_lpen       (rcc_c2_gpiog_lpen),
      .rcc_gpiof_arcg_clk_en   (rcc_gpiof_arcg_clk_en),
      .rcc_c1_gpiof_en         (rcc_c1_gpiof_en),
      .rcc_c2_gpiof_en         (rcc_c2_gpiof_en),
      .rcc_c1_gpiof_lpen       (rcc_c1_gpiof_lpen),
      .rcc_c2_gpiof_lpen       (rcc_c2_gpiof_lpen),
      .rcc_gpioe_arcg_clk_en   (rcc_gpioe_arcg_clk_en),
      .rcc_c1_gpioe_en         (rcc_c1_gpioe_en),
      .rcc_c2_gpioe_en         (rcc_c2_gpioe_en),
      .rcc_c1_gpioe_lpen       (rcc_c1_gpioe_lpen),
      .rcc_c2_gpioe_lpen       (rcc_c2_gpioe_lpen),
      .rcc_gpiod_arcg_clk_en   (rcc_gpiod_arcg_clk_en),
      .rcc_c1_gpiod_en         (rcc_c1_gpiod_en),
      .rcc_c2_gpiod_en         (rcc_c2_gpiod_en),
      .rcc_c1_gpiod_lpen       (rcc_c1_gpiod_lpen),
      .rcc_c2_gpiod_lpen       (rcc_c2_gpiod_lpen),
      .rcc_gpioc_arcg_clk_en   (rcc_gpioc_arcg_clk_en),
      .rcc_c1_gpioc_en         (rcc_c1_gpioc_en),
      .rcc_c2_gpioc_en         (rcc_c2_gpioc_en),
      .rcc_c1_gpioc_lpen       (rcc_c1_gpioc_lpen),
      .rcc_c2_gpioc_lpen       (rcc_c2_gpioc_lpen),
      .rcc_gpiob_arcg_clk_en   (rcc_gpiob_arcg_clk_en),
      .rcc_c1_gpiob_en         (rcc_c1_gpiob_en),
      .rcc_c2_gpiob_en         (rcc_c2_gpiob_en),
      .rcc_c1_gpiob_lpen       (rcc_c1_gpiob_lpen),
      .rcc_c2_gpiob_lpen       (rcc_c2_gpiob_lpen),
      .rcc_gpioa_arcg_clk_en   (rcc_gpioa_arcg_clk_en),
      .rcc_c1_gpioa_en         (rcc_c1_gpioa_en),
      .rcc_c2_gpioa_en         (rcc_c2_gpioa_en),
      .rcc_c1_gpioa_lpen       (rcc_c1_gpioa_lpen),
      .rcc_c2_gpioa_lpen       (rcc_c2_gpioa_lpen),
      .rcc_rcc_arcg_clk_en     (rcc_rcc_arcg_clk_en),
      .rcc_pwr_arcg_clk_en     (rcc_pwr_arcg_clk_en),
      .rcc_sai4_arcg_clk_en    (rcc_sai4_arcg_clk_en),
      .rcc_c1_sai4_en          (rcc_c1_sai4_en),
      .rcc_c2_sai4_en          (rcc_c2_sai4_en),
      .rcc_c1_sai4_lpen        (rcc_c1_sai4_lpen),
      .rcc_c2_sai4_lpen        (rcc_c2_sai4_lpen),
      .rcc_sai4_amen           (rcc_sai4_amen),
      .rcc_rtc_arcg_clk_en     (rcc_rtc_arcg_clk_en),
      .rcc_c1_rtc_en           (rcc_c1_rtc_en),
      .rcc_c2_rtc_en           (rcc_c2_rtc_en),
      .rcc_c1_rtc_lpen         (rcc_c1_rtc_lpen),
      .rcc_c2_rtc_lpen         (rcc_c2_rtc_lpen),
      .rcc_rtc_amen            (rcc_rtc_amen),
      .rcc_vref_arcg_clk_en    (rcc_vref_arcg_clk_en),
      .rcc_c1_vref_en          (rcc_c1_vref_en),
      .rcc_c2_vref_en          (rcc_c2_vref_en),
      .rcc_c1_vref_lpen        (rcc_c1_vref_lpen),
      .rcc_c2_vref_lpen        (rcc_c2_vref_lpen),
      .rcc_vref_amen           (rcc_vref_amen),
      .rcc_comp12_arcg_clk_en  (rcc_comp12_arcg_clk_en),
      .rcc_c1_comp12_en        (rcc_c1_comp12_en),
      .rcc_c2_comp12_en        (rcc_c2_comp12_en),
      .rcc_c1_comp12_lpen      (rcc_c1_comp12_lpen),
      .rcc_c2_comp12_lpen      (rcc_c2_comp12_lpen),
      .rcc_comp12_amen         (rcc_comp12_amen),
      .rcc_lptim5_arcg_clk_en  (rcc_lptim5_arcg_clk_en),
      .rcc_c1_lptim5_en        (rcc_c1_lptim5_en),
      .rcc_c2_lptim5_en        (rcc_c2_lptim5_en),
      .rcc_c1_lptim5_lpen      (rcc_c1_lptim5_lpen),
      .rcc_c2_lptim5_lpen      (rcc_c2_lptim5_lpen),
      .rcc_lptim5_amen         (rcc_lptim5_amen),
      .rcc_lptim4_arcg_clk_en  (rcc_lptim4_arcg_clk_en),
      .rcc_c1_lptim4_en        (rcc_c1_lptim4_en),
      .rcc_c2_lptim4_en        (rcc_c2_lptim4_en),
      .rcc_c1_lptim4_lpen      (rcc_c1_lptim4_lpen),
      .rcc_c2_lptim4_lpen      (rcc_c2_lptim4_lpen),
      .rcc_lptim4_amen         (rcc_lptim4_amen),
      .rcc_lptim3_arcg_clk_en  (rcc_lptim3_arcg_clk_en),
      .rcc_c1_lptim3_en        (rcc_c1_lptim3_en),
      .rcc_c2_lptim3_en        (rcc_c2_lptim3_en),
      .rcc_c1_lptim3_lpen      (rcc_c1_lptim3_lpen),
      .rcc_c2_lptim3_lpen      (rcc_c2_lptim3_lpen),
      .rcc_lptim3_amen         (rcc_lptim3_amen),
      .rcc_lptim2_arcg_clk_en  (rcc_lptim2_arcg_clk_en),
      .rcc_c1_lptim2_en        (rcc_c1_lptim2_en),
      .rcc_c2_lptim2_en        (rcc_c2_lptim2_en),
      .rcc_c1_lptim2_lpen      (rcc_c1_lptim2_lpen),
      .rcc_c2_lptim2_lpen      (rcc_c2_lptim2_lpen),
      .rcc_lptim2_amen         (rcc_lptim2_amen),
      .rcc_i2c4_arcg_clk_en    (rcc_i2c4_arcg_clk_en),
      .rcc_c1_i2c4_en          (rcc_c1_i2c4_en),
      .rcc_c2_i2c4_en          (rcc_c2_i2c4_en),
      .rcc_c1_i2c4_lpen        (rcc_c1_i2c4_lpen),
      .rcc_c2_i2c4_lpen        (rcc_c2_i2c4_lpen),
      .rcc_i2c4_amen           (rcc_i2c4_amen),
      .i2c4_ker_clk_req        (i2c4_ker_clk_req),
      .rcc_spi6_arcg_clk_en    (rcc_spi6_arcg_clk_en),
      .rcc_c1_spi6_en          (rcc_c1_spi6_en),
      .rcc_c2_spi6_en          (rcc_c2_spi6_en),
      .rcc_c1_spi6_lpen        (rcc_c1_spi6_lpen),
      .rcc_c2_spi6_lpen        (rcc_c2_spi6_lpen),
      .rcc_spi6_amen           (rcc_spi6_amen),
      .rcc_lpuart1_arcg_clk_en (rcc_lpuart1_arcg_clk_en),
      .rcc_c1_lpuart1_en       (rcc_c1_lpuart1_en),
      .rcc_c2_lpuart1_en       (rcc_c2_lpuart1_en),
      .rcc_c1_lpuart1_lpen     (rcc_c1_lpuart1_lpen),
      .rcc_c2_lpuart1_lpen     (rcc_c2_lpuart1_lpen),
      .rcc_lpuart1_amen        (rcc_lpuart1_amen),
      .lpuart1_ker_clk_req     (lpuart1_ker_clk_req),
      .rcc_syscfg_arcg_clk_en  (rcc_syscfg_arcg_clk_en),
      .rcc_c1_syscfg_en        (rcc_c1_syscfg_en),
      .rcc_c2_syscfg_en        (rcc_c2_syscfg_en),
      .rcc_c1_syscfg_lpen      (rcc_c1_syscfg_lpen),
      .rcc_c2_syscfg_lpen      (rcc_c2_syscfg_lpen),
      .rcc_iwdg2_arcg_clk_en   (rcc_iwdg2_arcg_clk_en),
      .rcc_iwdg1_arcg_clk_en   (rcc_iwdg1_arcg_clk_en),
      .rcc_exti_arcg_clk_en    (rcc_exti_arcg_clk_en),
      .qspisel                 (qspisel),
      .fmcsel                  (fmcsel),
      .sdmmcsel                (sdmmcsel),
      .usbsel                  (usbsel),
      .adcsel                  (adcsel),
      .rngsel                  (rngsel),
      .cecsel                  (cecsel),
      .i2c123sel               (i2c123sel),
      .usart234578sel          (usart234578sel),
      .spdifsel                (spdifsel),
      .lptim1sel               (lptim1sel),
      .fdcansel                (fdcansel),
      .swpmisel                (swpmisel),
      .sai1sel                 (sai1sel),
      .dfsdm1sel               (dfsdm1sel),
      .sai23sel                (sai23sel),
      .spi45sel                (spi45sel),
      .spi123sel               (spi123sel),
      .usart16sel              (usart16sel),
      .sai4asel                (sai4asel),
      .sai4bsel                (sai4bsel),
      .lptim345sel             (lptim345sel),
      .lptim2sel               (lptim2sel),
      .i2c4sel                 (i2c4sel),
      .spi6sel                 (spi6sel),
      .lpuart1sel              (lpuart1sel),

      .c2_per_alloc_d1     (c2_per_alloc_d1),
      .c1_per_alloc_d2     (c1_per_alloc_d2),
      .hsi_ker_clk_req     (hsi_ker_clk_req),
      .csi_ker_clk_req     (csi_ker_clk_req),
      .rcc_flash_aclk      (rcc_flash_aclk),
      .rcc_flash_hclk      (rcc_flash_hclk),
      .rcc_qspi_aclk       (rcc_qspi_aclk),
      .rcc_qspi_hclk       (rcc_qspi_hclk),
      .rcc_qspi_ker_clk    (rcc_qspi_ker_clk),
      .rcc_axisram_aclk    (rcc_axisram_aclk),
      .rcc_fmc_aclk        (rcc_fmc_aclk),
      .rcc_fmc_hclk        (rcc_fmc_hclk),
      .rcc_fmc_ker_clk     (rcc_fmc_ker_clk),
      .rcc_dma2d_aclk      (rcc_dma2d_aclk),
      .rcc_dma2d_hclk      (rcc_dma2d_hclk),
      .rcc_mdma_aclk       (rcc_mdma_aclk),
      .rcc_mdma_hclk       (rcc_mdma_hclk),
      .rcc_ltdc_aclk       (rcc_ltdc_aclk),
      .rcc_ltdc_pclk       (rcc_ltdc_pclk),
      .rcc_ltdc_ker_clk    (rcc_ltdc_ker_clk),
      .rcc_ramecc1_hclk    (rcc_ramecc1_hclk),
      .rcc_gpv_hclk        (rcc_gpv_hclk),
      .rcc_itcm_hclk       (rcc_itcm_hclk),
      .rcc_dtcm2_hclk      (rcc_dtcm2_hclk),
      .rcc_dtcm1_hclk      (rcc_dtcm1_hclk),
      .rcc_jpgdec_hclk     (rcc_jpgdec_hclk),
      .rcc_sdmmc1_hclk     (rcc_sdmmc1_hclk),
      .rcc_sdmmc1_ker_clk  (rcc_sdmmc1_ker_clk),
      .rcc_wwdg1_pclk      (rcc_wwdg1_pclk),
      .rcc_usb2ulpi_hclk   (rcc_usb2ulpi_hclk),
      .rcc_usb2otg_hclk    (rcc_usb2otg_hclk),
      .rcc_usb2otg_ker_clk (rcc_usb2otg_ker_clk),
      .rcc_usb1ulpi_hclk   (rcc_usb1ulpi_hclk),
      .rcc_usb1ulpi_ker_clk(rcc_usb1ulpi_ker_clk),
      .rcc_usb1otg_hclk    (rcc_usb1otg_hclk),
      .rcc_usb1otg_ker_clk (rcc_usb1otg_ker_clk),
      .rcc_eth1rx_hclk     (rcc_eth1rx_hclk),
      .rcc_eth1tx_hclk     (rcc_eth1tx_hclk),
      .rcc_eth1mac_hclk    (rcc_eth1mac_hclk),
      .rcc_adc12_hclk      (rcc_adc12_hclk),
      .rcc_adc12_ker_clk   (rcc_adc12_ker_clk),
      .rcc_dma2_hclk       (rcc_dma2_hclk),
      .rcc_dma1_hclk       (rcc_dma1_hclk),
      .rcc_sram3_hclk      (rcc_sram3_hclk),
      .rcc_sram2_hclk      (rcc_sram2_hclk),
      .rcc_sram1_hclk      (rcc_sram1_hclk),
      .rcc_sdmmc2_hclk     (rcc_sdmmc2_hclk),
      .rcc_sdmmc2_ker_clk  (rcc_sdmmc2_ker_clk),
      .rcc_rng_hclk        (rcc_rng_hclk),
      .rcc_rng_ker_clk     (rcc_rng_ker_clk),
      .rcc_hash_hclk       (rcc_hash_hclk),
      .rcc_crypt_hclk      (rcc_crypt_hclk),
      .rcc_dcmi_hclk       (rcc_dcmi_hclk),
      .rcc_ramecc2_hclk    (rcc_ramecc2_hclk),
      .rcc_uart8_pclk      (rcc_uart8_pclk),
      .rcc_uart8_ker_clk   (rcc_uart8_ker_clk),
      .rcc_uart7_pclk      (rcc_uart7_pclk),
      .rcc_uart7_ker_clk   (rcc_uart7_ker_clk),
      .rcc_dac12_pclk      (rcc_dac12_pclk),
      .rcc_hdmicec_pclk    (rcc_hdmicec_pclk),
      .rcc_hdmicec_ker_clk (rcc_hdmicec_ker_clk),
      .rcc_i2c3_pclk       (rcc_i2c3_pclk),
      .rcc_i2c3_ker_clk    (rcc_i2c3_ker_clk),
      .rcc_i2c2_pclk       (rcc_i2c2_pclk),
      .rcc_i2c2_ker_clk    (rcc_i2c2_ker_clk),
      .rcc_i2c1_pclk       (rcc_i2c1_pclk),
      .rcc_i2c1_ker_clk    (rcc_i2c1_ker_clk),
      .rcc_uart5_pclk      (rcc_uart5_pclk),
      .rcc_uart5_ker_clk   (rcc_uart5_ker_clk),
      .rcc_uart4_pclk      (rcc_uart4_pclk),
      .rcc_uart4_ker_clk   (rcc_uart4_ker_clk),
      .rcc_usart3_pclk     (rcc_usart3_pclk),
      .rcc_usart3_ker_clk  (rcc_usart3_ker_clk),
      .rcc_usart2_pclk     (rcc_usart2_pclk),
      .rcc_usart2_ker_clk  (rcc_usart2_ker_clk),
      .rcc_spdifrx_pclk    (rcc_spdifrx_pclk),
      .rcc_spdifrx_ker_clk (rcc_spdifrx_ker_clk),
      .rcc_spi3_pclk       (rcc_spi3_pclk),
      .rcc_spi3_ker_clk    (rcc_spi3_ker_clk),
      .rcc_spi2_pclk       (rcc_spi2_pclk),
      .rcc_spi2_ker_clk    (rcc_spi2_ker_clk),
      .rcc_wwdg2_pclk      (rcc_wwdg2_pclk),
      .rcc_lptim1_pclk     (rcc_lptim1_pclk),
      .rcc_lptim1_ker_clk  (rcc_lptim1_ker_clk),
      .rcc_tim14_pclk      (rcc_tim14_pclk),
      .rcc_tim14_ker_clk   (rcc_tim14_ker_clk),
      .rcc_tim13_pclk      (rcc_tim13_pclk),
      .rcc_tim13_ker_clk   (rcc_tim13_ker_clk),
      .rcc_tim12_pclk      (rcc_tim12_pclk),
      .rcc_tim12_ker_clk   (rcc_tim12_ker_clk),
      .rcc_tim7_pclk       (rcc_tim7_pclk),
      .rcc_tim7_ker_clk    (rcc_tim7_ker_clk),
      .rcc_tim6_pclk       (rcc_tim6_pclk),
      .rcc_tim6_ker_clk    (rcc_tim6_ker_clk),
      .rcc_tim5_pclk       (rcc_tim5_pclk),
      .rcc_tim5_ker_clk    (rcc_tim5_ker_clk),
      .rcc_tim4_pclk       (rcc_tim4_pclk),
      .rcc_tim4_ker_clk    (rcc_tim4_ker_clk),
      .rcc_tim3_pclk       (rcc_tim3_pclk),
      .rcc_tim3_ker_clk    (rcc_tim3_ker_clk),
      .rcc_tim2_pclk       (rcc_tim2_pclk),
      .rcc_tim2_ker_clk    (rcc_tim2_ker_clk),
      .rcc_fdcan_pclk      (rcc_fdcan_pclk),
      .rcc_fdcan_ker_clk   (rcc_fdcan_ker_clk),
      .rcc_mdios_pclk      (rcc_mdios_pclk),
      .rcc_opamp_pclk      (rcc_opamp_pclk),
      .rcc_swpmi_pclk      (rcc_swpmi_pclk),
      .rcc_swpmi_ker_clk   (rcc_swpmi_ker_clk),
      .rcc_crs_pclk        (rcc_crs_pclk),
      .rcc_hrtim_pclk      (rcc_hrtim_pclk),
      .rcc_hrtim_ker_clk   (rcc_hrtim_ker_clk),
      .rcc_dfsdm1_pclk     (rcc_dfsdm1_pclk),
      .rcc_dfsdm1_ker_clk_0(rcc_dfsdm1_ker_clk_0),
      .rcc_dfsdm1_ker_clk_1(rcc_dfsdm1_ker_clk_1),
      .rcc_sai3_pclk       (rcc_sai3_pclk),
      .rcc_sai3_ker_clk    (rcc_sai3_ker_clk),
      .rcc_sai2_pclk       (rcc_sai2_pclk),
      .rcc_sai2_ker_clk    (rcc_sai2_ker_clk),
      .rcc_sai1_pclk       (rcc_sai1_pclk),
      .rcc_sai1_ker_clk    (rcc_sai1_ker_clk),
      .rcc_spi5_pclk       (rcc_spi5_pclk),
      .rcc_spi5_ker_clk    (rcc_spi5_ker_clk),
      .rcc_tim17_pclk      (rcc_tim17_pclk),
      .rcc_tim17_ker_clk   (rcc_tim17_ker_clk),
      .rcc_tim16_pclk      (rcc_tim16_pclk),
      .rcc_tim16_ker_clk   (rcc_tim16_ker_clk),
      .rcc_tim15_pclk      (rcc_tim15_pclk),
      .rcc_tim15_ker_clk   (rcc_tim15_ker_clk),
      .rcc_spi4_pclk       (rcc_spi4_pclk),
      .rcc_spi4_ker_clk    (rcc_spi4_ker_clk),
      .rcc_spi1_pclk       (rcc_spi1_pclk),
      .rcc_spi1_ker_clk    (rcc_spi1_ker_clk),
      .rcc_usart6_pclk     (rcc_usart6_pclk),
      .rcc_usart6_ker_clk  (rcc_usart6_ker_clk),
      .rcc_usart1_pclk     (rcc_usart1_pclk),
      .rcc_usart1_ker_clk  (rcc_usart1_ker_clk),
      .rcc_tim8_pclk       (rcc_tim8_pclk),
      .rcc_tim8_ker_clk    (rcc_tim8_ker_clk),
      .rcc_tim1_pclk       (rcc_tim1_pclk),
      .rcc_tim1_ker_clk    (rcc_tim1_ker_clk),
      .rcc_sram4_hclk      (rcc_sram4_hclk),
      .rcc_bkpram_hclk     (rcc_bkpram_hclk),
      .rcc_ramecc3_hclk    (rcc_ramecc3_hclk),
      .rcc_hsem_hclk       (rcc_hsem_hclk),
      .rcc_adc3_hclk       (rcc_adc3_hclk),
      .rcc_adc3_ker_clk    (rcc_adc3_ker_clk),
      .rcc_bdma_hclk       (rcc_bdma_hclk),
      .rcc_crc_hclk        (rcc_crc_hclk),
      .rcc_gpiok_hclk      (rcc_gpiok_hclk),
      .rcc_gpioj_hclk      (rcc_gpioj_hclk),
      .rcc_gpioi_hclk      (rcc_gpioi_hclk),
      .rcc_gpioh_hclk      (rcc_gpioh_hclk),
      .rcc_gpiog_hclk      (rcc_gpiog_hclk),
      .rcc_gpiof_hclk      (rcc_gpiof_hclk),
      .rcc_gpioe_hclk      (rcc_gpioe_hclk),
      .rcc_gpiod_hclk      (rcc_gpiod_hclk),
      .rcc_gpioc_hclk      (rcc_gpioc_hclk),
      .rcc_gpiob_hclk      (rcc_gpiob_hclk),
      .rcc_gpioa_hclk      (rcc_gpioa_hclk),
      .rcc_rcc_hclk        (rcc_rcc_hclk),
      .rcc_pwr_hclk        (rcc_pwr_hclk),
      .rcc_sai4_pclk       (rcc_sai4_pclk),
      .rcc_sai4_ker_clk_0  (rcc_sai4_ker_clk_0),
      .rcc_sai4_ker_clk_1  (rcc_sai4_ker_clk_1),
      .rcc_rtc_pclk        (rcc_rtc_pclk),
      .rcc_vref_pclk       (rcc_vref_pclk),
      .rcc_comp12_pclk     (rcc_comp12_pclk),
      .rcc_lptim5_pclk     (rcc_lptim5_pclk),
      .rcc_lptim5_ker_clk  (rcc_lptim5_ker_clk),
      .rcc_lptim4_pclk     (rcc_lptim4_pclk),
      .rcc_lptim4_ker_clk  (rcc_lptim4_ker_clk),
      .rcc_lptim3_pclk     (rcc_lptim3_pclk),
      .rcc_lptim3_ker_clk  (rcc_lptim3_ker_clk),
      .rcc_lptim2_pclk     (rcc_lptim2_pclk),
      .rcc_lptim2_ker_clk  (rcc_lptim2_ker_clk),
      .rcc_i2c4_pclk       (rcc_i2c4_pclk),
      .rcc_i2c4_ker_clk    (rcc_i2c4_ker_clk),
      .rcc_spi6_pclk       (rcc_spi6_pclk),
      .rcc_spi6_ker_clk    (rcc_spi6_ker_clk),
      .rcc_lpuart1_pclk    (rcc_lpuart1_pclk),
      .rcc_lpuart1_ker_clk (rcc_lpuart1_ker_clk),
      .rcc_syscfg_pclk     (rcc_syscfg_pclk),
      .rcc_iwdg2_pclk      (rcc_iwdg2_pclk),
      .rcc_iwdg1_pclk      (rcc_iwdg1_pclk),
      .rcc_exti_pclk       (rcc_exti_pclk)
  );


endmodule
