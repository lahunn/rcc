module rcc_top #(
    parameter CLK_ON_AFTER_PER_RST_RELEASE  = 8,
    parameter CLK_ON_AFTER_SYS_RST_RELEASE  = 8,
    parameter CLK_ON_AFTER_D1_RST_RELEASE   = 8,
    parameter CLK_ON_AFTER_D2_RST_RELEASE   = 8,
    parameter CLK_ON_AFTER_CPU1_RST_RELEASE = 8,
    parameter CLK_ON_AFTER_CPU2_RST_RELEASE = 8
) (
    // signals connected to 复位源 
    input  nrst_in,
    input  iwdg1_out_rst,
    input  wwdg1_out_rst,
    input  iwdg2_out_rst,
    input  wwdg2_out_rst,
    input  lpwr2_rst,
    input  lpwr1_rst,
    input  pwr_bor_rst,
    input  pwr_por_rst,
    input  cpu2_sftrst,
    input  cpu1_sftrst,
    output nrst_out,

    // signals connected to PWR 
    input  d3_deepsleep,
    input  pwr_d1_wkup,
    input  pwr_d2_wkup,
    input  pwr_d3_wkup,
    output rcc_pwr_d1_req,
    output rcc_pwr_d2_req,
    output rcc_pwr_d3_req,
    output c2_per_alloc_d1,
    output c1_per_alloc_d2,
    input  flash_power_ok,
    input  pwr_d1_ok,
    input  pwr_d2_ok,
    input  pwr_vcore_ok,
    input  backup_protect,


    // signals connected to CPU 
    input  c2_sleep,
    input  c2_deepsleep,
    input  c1_sleep,
    input  c1_deepsleep,
    output rcc_c2_clk,
    output rcc_fclk_c2,
    output rcc_c2_systick_clk,
    output rcc_c1_clk,
    output rcc_fclk_c1,
    output rcc_c1_systick_clk,
    // reset to cpu and bus 
    output cpu1_arcg_rst_n,
    output cpu2_arcg_rst_n,
    output d1_bus_arcg_rst_n,
    output d2_bus_arcg_rst_n,
    output d3_bus_arcg_rst_n,
    // timer clocks
    output rcc_timx_ker_clk,
    output rcc_timy_ker_clk,
    output rcc_hrtimer_prescalar_clk,
    output sys_d1cpre_clk,
    output sys_hpre_clk,
    // signals connected to PAD 
    output mco1,
    output mco2,
    input  pad_rcc_eth_mii_tx_clk,
    input  pad_rcc_eth_mii_rx_clk,
    input  USB_PHY1,
    // interrupt signals
    output rcc_hsefail_it,
    output rcc_lsefail_it,
    output rcc_it,

    // some other signals 
    input        flash_obl_reload,
    input        obl_done,
    input        rcc_arcg_on,
    input        pll3_rdy,
    input        pll2_rdy,
    input        pll1_rdy,
    input        hse_rdy,
    input        hsi48_rdy,
    input        csi_rdy,
    input        hsi_rdy,
    input [ 7:0] flash_csi_opt,
    input [11:0] flash_hsi_opt,
    input [ 9:0] crs_hsi48_trim,
    input        rcc_hsecss_fail,
    input        rcc_lsecss_fail,


    // reset signals
    output pwr_por_rst_n,
    output sys_arcg_rst_n,
    output d1_arcg_rst_n,
    output d2_arcg_rst_n,
    output stby_rst_n,

    // per rst signals
    output        rcc_flash_arcg_rst_n,
    output        rcc_qspi_arcg_rst_n,
    output        rcc_axisram_arcg_rst_n,
    output        rcc_fmc_arcg_rst_n,
    output        rcc_dma2d_arcg_rst_n,
    output        rcc_mdma_arcg_rst_n,
    output        rcc_ltdc_arcg_rst_n,
    output        rcc_ramecc1_arcg_rst_n,
    output        rcc_gpv_arcg_rst_n,
    output        rcc_itcm_arcg_rst_n,
    output        rcc_dtcm2_arcg_rst_n,
    output        rcc_dtcm1_arcg_rst_n,
    output        rcc_jpgdec_arcg_rst_n,
    output        rcc_sdmmc1_arcg_rst_n,
    output        rcc_wwdg1_arcg_rst_n,
    output        rcc_usb2ulpi_arcg_rst_n,
    output        rcc_usb2otg_arcg_rst_n,
    output        rcc_usb1ulpi_arcg_rst_n,
    output        rcc_usb1otg_arcg_rst_n,
    output        rcc_eth1rx_arcg_rst_n,
    output        rcc_eth1tx_arcg_rst_n,
    output        rcc_eth1mac_arcg_rst_n,
    output        rcc_adc12_arcg_rst_n,
    output        rcc_dma2_arcg_rst_n,
    output        rcc_dma1_arcg_rst_n,
    output        rcc_sram3_arcg_rst_n,
    output        rcc_sram2_arcg_rst_n,
    output        rcc_sram1_arcg_rst_n,
    output        rcc_sdmmc2_arcg_rst_n,
    output        rcc_rng_arcg_rst_n,
    output        rcc_hash_arcg_rst_n,
    output        rcc_crypt_arcg_rst_n,
    output        rcc_dcmi_arcg_rst_n,
    output        rcc_ramecc2_arcg_rst_n,
    output        rcc_uart8_arcg_rst_n,
    output        rcc_uart7_arcg_rst_n,
    output        rcc_dac12_arcg_rst_n,
    output        rcc_hdmicec_arcg_rst_n,
    output        rcc_i2c3_arcg_rst_n,
    output        rcc_i2c2_arcg_rst_n,
    output        rcc_i2c1_arcg_rst_n,
    output        rcc_uart5_arcg_rst_n,
    output        rcc_uart4_arcg_rst_n,
    output        rcc_usart3_arcg_rst_n,
    output        rcc_usart2_arcg_rst_n,
    output        rcc_spdifrx_arcg_rst_n,
    output        rcc_spi3_arcg_rst_n,
    output        rcc_spi2_arcg_rst_n,
    output        rcc_wwdg2_arcg_rst_n,
    output        rcc_lptim1_arcg_rst_n,
    output        rcc_tim14_arcg_rst_n,
    output        rcc_tim13_arcg_rst_n,
    output        rcc_tim12_arcg_rst_n,
    output        rcc_tim7_arcg_rst_n,
    output        rcc_tim6_arcg_rst_n,
    output        rcc_tim5_arcg_rst_n,
    output        rcc_tim4_arcg_rst_n,
    output        rcc_tim3_arcg_rst_n,
    output        rcc_tim2_arcg_rst_n,
    output        rcc_fdcan_arcg_rst_n,
    output        rcc_mdios_arcg_rst_n,
    output        rcc_opamp_arcg_rst_n,
    output        rcc_swpmi_arcg_rst_n,
    output        rcc_crs_arcg_rst_n,
    output        rcc_hrtim_arcg_rst_n,
    output        rcc_dfsdm1_arcg_rst_n,
    output        rcc_sai3_arcg_rst_n,
    output        rcc_sai2_arcg_rst_n,
    output        rcc_sai1_arcg_rst_n,
    output        rcc_spi5_arcg_rst_n,
    output        rcc_tim17_arcg_rst_n,
    output        rcc_tim16_arcg_rst_n,
    output        rcc_tim15_arcg_rst_n,
    output        rcc_spi4_arcg_rst_n,
    output        rcc_spi1_arcg_rst_n,
    output        rcc_usart6_arcg_rst_n,
    output        rcc_usart1_arcg_rst_n,
    output        rcc_tim8_arcg_rst_n,
    output        rcc_tim1_arcg_rst_n,
    output        rcc_sram4_arcg_rst_n,
    output        rcc_bkpram_arcg_rst_n,
    output        rcc_ramecc3_arcg_rst_n,
    output        rcc_hsem_arcg_rst_n,
    output        rcc_adc3_arcg_rst_n,
    output        rcc_bdma_arcg_rst_n,
    output        rcc_crc_arcg_rst_n,
    output        rcc_gpiok_arcg_rst_n,
    output        rcc_gpioj_arcg_rst_n,
    output        rcc_gpioi_arcg_rst_n,
    output        rcc_gpioh_arcg_rst_n,
    output        rcc_gpiog_arcg_rst_n,
    output        rcc_gpiof_arcg_rst_n,
    output        rcc_gpioe_arcg_rst_n,
    output        rcc_gpiod_arcg_rst_n,
    output        rcc_gpioc_arcg_rst_n,
    output        rcc_gpiob_arcg_rst_n,
    output        rcc_gpioa_arcg_rst_n,
    output        rcc_rcc_arcg_rst_n,
    output        rcc_pwr_arcg_rst_n,
    output        rcc_sai4_arcg_rst_n,
    output        rcc_rtc_arcg_rst_n,
    output        rcc_vref_arcg_rst_n,
    output        rcc_comp12_arcg_rst_n,
    output        rcc_lptim5_arcg_rst_n,
    output        rcc_lptim4_arcg_rst_n,
    output        rcc_lptim3_arcg_rst_n,
    output        rcc_lptim2_arcg_rst_n,
    output        rcc_i2c4_arcg_rst_n,
    output        rcc_spi6_arcg_rst_n,
    output        rcc_lpuart1_arcg_rst_n,
    output        rcc_syscfg_arcg_rst_n,
    output        rcc_iwdg2_arcg_rst_n,
    output        rcc_iwdg1_arcg_rst_n,
    output        rcc_exti_arcg_rst_n,
    // ahb bus signals
    input         ahb_hclk,
    input         ahb_hresetn,
    input  [31:0] ahb_haddr,
    input  [ 2:0] ahb_hburst,
    input  [ 2:0] ahb_hprot,
    output [31:0] ahb_hrdata,
    input         ahb_hready_in,
    output        ahb_hready_out,
    output        ahb_hresp,
    input  [ 2:0] ahb_hsize,
    input  [ 1:0] ahb_htrans,
    input  [31:0] ahb_hwdata,
    input         ahb_hwrite,
    input         ahb_hsel,
    input         ahb_hmaster,

    // per_ker_clk_control Inputs
    // ker clock req
    input         uart8_ker_clk_req,
    input         uart7_ker_clk_req,
    input         i2c3_ker_clk_req,
    input         i2c2_ker_clk_req,
    input         i2c1_ker_clk_req,
    input         uart5_ker_clk_req,
    input         uart4_ker_clk_req,
    input         usart3_ker_clk_req,
    input         usart2_ker_clk_req,
    input         usart6_ker_clk_req,
    input         usart1_ker_clk_req,
    input         i2c4_ker_clk_req,
    input         lpuart1_ker_clk_req,
    // bus clock signals
    output        rcc_axibridge_d1_clk,
    output        rcc_ahb3bridge_d1_clk,
    output        rcc_apb3bridge_d1_clk,
    output        rcc_ahb1bridge_d2_clk,
    output        rcc_ahb2bridge_d2_clk,
    output        rcc_apb1bridge_d2_clk,
    output        rcc_apb2bridge_d2_clk,
    output        rcc_ahb4bridge_d3_clk,
    output        rcc_apb4bridge_d3_clk,
    // pll , oscilator and pad clocks
    output        pll1_src_clk,
    output        pll2_src_clk,
    output        pll3_src_clk,
    input         pll1_p_clk,
    input         pll1_q_clk,
    input         pll2_p_clk,
    input         pll2_q_clk,
    input         pll2_r_clk,
    input         pll3_p_clk,
    input         pll3_q_clk,
    input         pll3_r_clk,
    input         I2S_clk_IN,
    // pll osc control signals
    output        pll3on,
    output        pll2on,
    output        pll1on,
    output        hsecsson,
    output        hsebyp,
    output        hseon,
    output        hsi48on,
    output        csikeron,
    output        csion,
    output [ 1:0] hsidiv,
    output        hsikeron,
    output        hsion,
    output [ 7:0] rcc_csi_triming,
    output [11:0] rcc_hsi_triming,
    output        divr3en,
    output        divq3en,
    output        divp3en,
    output        divr2en,
    output        divq2en,
    output        divp2en,
    output        divr1en,
    output        divq1en,
    output        divp1en,
    output [ 1:0] pll3rge,
    output        pll3vcosel,
    output        pll3fracen,
    output [ 1:0] pll2rge,
    output        pll2vcosel,
    output        pll2fracen,
    output [ 1:0] pll1rge,
    output        pll1vcosel,
    output        pll1fracen,
    output [ 6:0] divr1,
    output [ 6:0] divq1,
    output [ 6:0] divp1,
    output [ 8:0] divn1,
    output [12:0] fracn1,
    output [ 6:0] divr2,
    output [ 6:0] divq2,
    output [ 6:0] divp2,
    output [ 8:0] divn2,
    output [12:0] fracn2,
    output [ 6:0] divr3,
    output [ 6:0] divq3,
    output [ 6:0] divp3,
    output [ 8:0] divn3,
    output [12:0] fracn3,
    // indicate busy state 
    input         axibridge_d1_busy,
    input         ahb3bridge_d1_busy,
    input         apb3bridge_d1_busy,
    input         ahb1bridge_d2_busy,
    input         ahb2bridge_d2_busy,
    input         apb1bridge_d2_busy,
    input         apb2bridge_d2_busy,
    input         ahb4bridge_d3_busy,
    input         apb4bridge_d3_busy,
    input         flash_busy,
    // signals connected to HSE
    input         hse_css_fail,
    input         hse_clk_pre,
    // lse lsi clock
    input         lse_clk,
    input         lsi_clk,
    // signals connected to HSI48 
    input         hsi48_clk,
    // signals connected to CSI
    input         csi_clk_pre,
    // signals connected to HSI
    input         hsi_origin_clk,
    //signals from eth 
    input         eth_rcc_fes,
    input         eth_rcc_epis_2,
    output        rcc_eth_mii_tx_clk,
    output        rcc_eth_mii_rx_clk,
    output        rcc_eth_rmii_ref_clk,

    //per_ker_clk_control region
    output       rcc_rtc_pclk,
    output       rcc_flash_aclk,
    output       rcc_flash_hclk,
    output       rcc_qspi_aclk,
    output       rcc_qspi_hclk,
    output       rcc_qspi_ker_clk,
    output       rcc_axisram_aclk,
    output       rcc_fmc_aclk,
    output       rcc_fmc_hclk,
    output       rcc_fmc_ker_clk,
    output       rcc_dma2d_aclk,
    output       rcc_dma2d_hclk,
    output       rcc_mdma_aclk,
    output       rcc_mdma_hclk,
    output       rcc_ltdc_aclk,
    output       rcc_ltdc_pclk,
    output       rcc_ltdc_ker_clk,
    output       rcc_ramecc1_hclk,
    output       rcc_gpv_hclk,
    output       rcc_itcm_hclk,
    output       rcc_dtcm2_hclk,
    output       rcc_dtcm1_hclk,
    output       rcc_jpgdec_hclk,
    output       rcc_sdmmc1_hclk,
    output       rcc_sdmmc1_ker_clk,
    output       rcc_wwdg1_pclk,
    output       rcc_usb2ulpi_hclk,
    output       rcc_usb2otg_hclk,
    output       rcc_usb2otg_ker_clk,
    output       rcc_usb1ulpi_hclk,
    output       rcc_usb1ulpi_ker_clk,
    output       rcc_usb1otg_hclk,
    output       rcc_usb1otg_ker_clk,
    output       rcc_eth1rx_hclk,
    output       rcc_eth1tx_hclk,
    output       rcc_eth1mac_hclk,
    output       rcc_adc12_hclk,
    output       rcc_adc12_ker_clk,
    output       rcc_dma2_hclk,
    output       rcc_dma1_hclk,
    output       rcc_sram3_hclk,
    output       rcc_sram2_hclk,
    output       rcc_sram1_hclk,
    output       rcc_sdmmc2_hclk,
    output       rcc_sdmmc2_ker_clk,
    output       rcc_rng_hclk,
    output       rcc_rng_ker_clk,
    output       rcc_hash_hclk,
    output       rcc_crypt_hclk,
    output       rcc_dcmi_hclk,
    output       rcc_ramecc2_hclk,
    output       rcc_uart8_pclk,
    output       rcc_uart8_ker_clk,
    output       rcc_uart7_pclk,
    output       rcc_uart7_ker_clk,
    output       rcc_dac12_pclk,
    output       rcc_hdmicec_pclk,
    output       rcc_hdmicec_ker_clk,
    output       rcc_i2c3_pclk,
    output       rcc_i2c3_ker_clk,
    output       rcc_i2c2_pclk,
    output       rcc_i2c2_ker_clk,
    output       rcc_i2c1_pclk,
    output       rcc_i2c1_ker_clk,
    output       rcc_uart5_pclk,
    output       rcc_uart5_ker_clk,
    output       rcc_uart4_pclk,
    output       rcc_uart4_ker_clk,
    output       rcc_usart3_pclk,
    output       rcc_usart3_ker_clk,
    output       rcc_usart2_pclk,
    output       rcc_usart2_ker_clk,
    output       rcc_spdifrx_pclk,
    output       rcc_spdifrx_ker_clk,
    output       rcc_spi3_pclk,
    output       rcc_spi3_ker_clk,
    output       rcc_spi2_pclk,
    output       rcc_spi2_ker_clk,
    output       rcc_wwdg2_pclk,
    output       rcc_lptim1_pclk,
    output       rcc_lptim1_ker_clk,
    output       rcc_tim14_pclk,
    output       rcc_tim14_ker_clk,
    output       rcc_tim13_pclk,
    output       rcc_tim13_ker_clk,
    output       rcc_tim12_pclk,
    output       rcc_tim12_ker_clk,
    output       rcc_tim7_pclk,
    output       rcc_tim7_ker_clk,
    output       rcc_tim6_pclk,
    output       rcc_tim6_ker_clk,
    output       rcc_tim5_pclk,
    output       rcc_tim5_ker_clk,
    output       rcc_tim4_pclk,
    output       rcc_tim4_ker_clk,
    output       rcc_tim3_pclk,
    output       rcc_tim3_ker_clk,
    output       rcc_tim2_pclk,
    output       rcc_tim2_ker_clk,
    output       rcc_fdcan_pclk,
    output       rcc_fdcan_ker_clk,
    output       rcc_mdios_pclk,
    output       rcc_opamp_pclk,
    output       rcc_swpmi_pclk,
    output       rcc_swpmi_ker_clk,
    output       rcc_crs_pclk,
    output       rcc_hrtim_pclk,
    output       rcc_hrtim_ker_clk,
    output       rcc_dfsdm1_pclk,
    output       rcc_dfsdm1_ker_clk_0,
    output       rcc_dfsdm1_ker_clk_1,
    output       rcc_sai3_pclk,
    output       rcc_sai3_ker_clk,
    output       rcc_sai2_pclk,
    output       rcc_sai2_ker_clk,
    output       rcc_sai1_pclk,
    output       rcc_sai1_ker_clk,
    output       rcc_spi5_pclk,
    output       rcc_spi5_ker_clk,
    output       rcc_tim17_pclk,
    output       rcc_tim17_ker_clk,
    output       rcc_tim16_pclk,
    output       rcc_tim16_ker_clk,
    output       rcc_tim15_pclk,
    output       rcc_tim15_ker_clk,
    output       rcc_spi4_pclk,
    output       rcc_spi4_ker_clk,
    output       rcc_spi1_pclk,
    output       rcc_spi1_ker_clk,
    output       rcc_usart6_pclk,
    output       rcc_usart6_ker_clk,
    output       rcc_usart1_pclk,
    output       rcc_usart1_ker_clk,
    output       rcc_tim8_pclk,
    output       rcc_tim8_ker_clk,
    output       rcc_tim1_pclk,
    output       rcc_tim1_ker_clk,
    output       rcc_sram4_hclk,
    output       rcc_bkpram_hclk,
    output       rcc_ramecc3_hclk,
    output       rcc_hsem_hclk,
    output       rcc_adc3_hclk,
    output       rcc_adc3_ker_clk,
    output       rcc_bdma_hclk,
    output       rcc_crc_hclk,
    output       rcc_gpiok_hclk,
    output       rcc_gpioj_hclk,
    output       rcc_gpioi_hclk,
    output       rcc_gpioh_hclk,
    output       rcc_gpiog_hclk,
    output       rcc_gpiof_hclk,
    output       rcc_gpioe_hclk,
    output       rcc_gpiod_hclk,
    output       rcc_gpioc_hclk,
    output       rcc_gpiob_hclk,
    output       rcc_gpioa_hclk,
    output       rcc_rcc_hclk,
    output       rcc_pwr_hclk,
    output       rcc_sai4_pclk,
    output       rcc_sai4_ker_clk_0,
    output       rcc_sai4_ker_clk_1,
    output       rcc_vref_pclk,
    output       rcc_comp12_pclk,
    output       rcc_lptim5_pclk,
    output       rcc_lptim5_ker_clk,
    output       rcc_lptim4_pclk,
    output       rcc_lptim4_ker_clk,
    output       rcc_lptim3_pclk,
    output       rcc_lptim3_ker_clk,
    output       rcc_lptim2_pclk,
    output       rcc_lptim2_ker_clk,
    output       rcc_i2c4_pclk,
    output       rcc_i2c4_ker_clk,
    output       rcc_spi6_pclk,
    output       rcc_spi6_ker_clk,
    output       rcc_lpuart1_pclk,
    output       rcc_lpuart1_ker_clk,
    output       rcc_syscfg_pclk,
    output       rcc_iwdg2_pclk,
    output       rcc_iwdg1_pclk,
    output       rcc_exti_pclk,
    // lse signal 
    output       lsecss_fail,
    input        lserdy,
    input        pwr_vsw_rst,
    output       bdrst,
    output       rtcen,
    output [1:0] rtcsel,
    output       lsecssd,
    output       lsecsson,
    output [1:0] lsedrv,
    output       lsebyp,
    output       lseon
);

  // rcc_vsw_top Inputs
  wire       hse_rtc_clk;
  wire       rcc_bdcr_byte2_wren;
  wire       rcc_bdcr_byte1_wren;
  wire       rcc_bdcr_byte0_wren;
  wire       nxt_rcc_bdcr_bdrst;
  wire       nxt_rcc_bdcr_rtcen;
  wire [1:0] nxt_rcc_bdcr_rtcsel;
  wire       nxt_rcc_bdcr_lsecsson;
  wire [1:0] nxt_rcc_bdcr_lsedrv;
  wire       nxt_rcc_bdcr_lsebyp;
  wire       nxt_rcc_bdcr_lseon;

  // rcc_vsw_top Outputs
  wire       rcc_rtc_ker_clk;
  wire       cur_rcc_bdcr_lserdy;

  // rcc_vdd_top Inputs
  wire       vdd_wdata;
  wire       rcc_c1_rsr_rmvf_wren;
  wire       rcc_c2_rsr_rmvf_wren;
  wire       rcc_csr_lsion_wren;
  wire       obl_rst;

  wire       d2_rst;
  wire       d1_rst;
  wire       lsi_rdy;

  // rcc_vdd_top Outputs
  wire       cur_rcc_c1_rsr_lpwr2rstf;
  wire       cur_rcc_c1_rsr_lpwr1rstf;
  wire       cur_rcc_c1_rsr_wwdg2rstf;
  wire       cur_rcc_c1_rsr_wwdg1rstf;
  wire       cur_rcc_c1_rsr_iwdg2rstf;
  wire       cur_rcc_c1_rsr_iwdg1rstf;
  wire       cur_rcc_c1_rsr_sft2rstf;
  wire       cur_rcc_c1_rsr_sft1rstf;
  wire       cur_rcc_c1_rsr_porrstf;
  wire       cur_rcc_c1_rsr_pinrstf;
  wire       cur_rcc_c1_rsr_borrstf;
  wire       cur_rcc_c1_rsr_d2rstf;
  wire       cur_rcc_c1_rsr_d1rstf;
  wire       cur_rcc_c1_rsr_oblrstf;
  wire       cur_rcc_c1_rsr_rmvf;
  wire       cur_rcc_c2_rsr_lpwr2rstf;
  wire       cur_rcc_c2_rsr_lpwr1rstf;
  wire       cur_rcc_c2_rsr_wwdg2rstf;
  wire       cur_rcc_c2_rsr_wwdg1rstf;
  wire       cur_rcc_c2_rsr_iwdg2rstf;
  wire       cur_rcc_c2_rsr_iwdg1rstf;
  wire       cur_rcc_c2_rsr_sft2rstf;
  wire       cur_rcc_c2_rsr_sft1rstf;
  wire       cur_rcc_c2_rsr_porrstf;
  wire       cur_rcc_c2_rsr_pinrstf;
  wire       cur_rcc_c2_rsr_borrstf;
  wire       cur_rcc_c2_rsr_d2rstf;
  wire       cur_rcc_c2_rsr_d1rstf;
  wire       cur_rcc_c2_rsr_oblrstf;
  wire       cur_rcc_c2_rsr_rmvf;
  wire       cur_rcc_csr_lsirdy;
  wire       cur_rcc_csr_lsion;

  rcc_vsw_top u_rcc_vsw_top (
      .lsecss_fail          (lsecss_fail),
      .lse_clk              (lse_clk),
      .lserdy               (lserdy),
      .lsi_clk              (lsi_clk),
      .hse_rtc_clk          (hse_rtc_clk),
      .pwr_vsw_rst          (pwr_vsw_rst),
      .rcc_bdcr_byte2_wren  (rcc_bdcr_byte2_wren),
      .rcc_bdcr_byte1_wren  (rcc_bdcr_byte1_wren),
      .rcc_bdcr_byte0_wren  (rcc_bdcr_byte0_wren),
      .nxt_rcc_bdcr_bdrst   (nxt_rcc_bdcr_bdrst),
      .nxt_rcc_bdcr_rtcen   (nxt_rcc_bdcr_rtcen),
      .nxt_rcc_bdcr_rtcsel  (nxt_rcc_bdcr_rtcsel),
      .nxt_rcc_bdcr_lsecsson(nxt_rcc_bdcr_lsecsson),
      .nxt_rcc_bdcr_lsedrv  (nxt_rcc_bdcr_lsedrv),
      .nxt_rcc_bdcr_lsebyp  (nxt_rcc_bdcr_lsebyp),
      .nxt_rcc_bdcr_lseon   (nxt_rcc_bdcr_lseon),

      .rcc_rtc_ker_clk    (rcc_rtc_ker_clk),
      .bdrst              (bdrst),
      .rtcen              (rtcen),
      .rtcsel             (rtcsel),
      .lsecssd            (lsecssd),
      .lsecsson           (lsecsson),
      .lsedrv             (lsedrv),
      .lsebyp             (lsebyp),
      .cur_rcc_bdcr_lserdy(cur_rcc_bdcr_lserdy),
      .lseon              (lseon)
  );

  rcc_vdd_top u_rcc_vdd_top (
      .wdata               (wdata),
      .rcc_c1_rsr_rmvf_wren(rcc_c1_rsr_rmvf_wren),
      .rcc_c2_rsr_rmvf_wren(rcc_c2_rsr_rmvf_wren),
      .rcc_csr_lsion_wren  (rcc_csr_lsion_wren),
      .nrst_in             (nrst_in),
      .obl_rst             (obl_rst),
      .lpwr2_rst           (lpwr2_rst),
      .lpwr1_rst           (lpwr1_rst),
      .wwdg1_out_rst       (wwdg1_out_rst),
      .wwdg2_out_rst       (wwdg2_out_rst),
      .iwdg1_out_rst       (iwdg1_out_rst),
      .iwdg2_out_rst       (iwdg2_out_rst),
      .cpu2_sftrst         (cpu2_sftrst),
      .cpu1_sftrst         (cpu1_sftrst),
      .pwr_por_rst         (pwr_por_rst),
      .pwr_bor_rst         (pwr_bor_rst),
      .d2_rst              (d2_rst),
      .d1_rst              (d1_rst),
      .lsi_rdy             (lsi_rdy),

      .cur_rcc_c1_rsr_lpwr2rstf(cur_rcc_c1_rsr_lpwr2rstf),
      .cur_rcc_c1_rsr_lpwr1rstf(cur_rcc_c1_rsr_lpwr1rstf),
      .cur_rcc_c1_rsr_wwdg2rstf(cur_rcc_c1_rsr_wwdg2rstf),
      .cur_rcc_c1_rsr_wwdg1rstf(cur_rcc_c1_rsr_wwdg1rstf),
      .cur_rcc_c1_rsr_iwdg2rstf(cur_rcc_c1_rsr_iwdg2rstf),
      .cur_rcc_c1_rsr_iwdg1rstf(cur_rcc_c1_rsr_iwdg1rstf),
      .cur_rcc_c1_rsr_sft2rstf (cur_rcc_c1_rsr_sft2rstf),
      .cur_rcc_c1_rsr_sft1rstf (cur_rcc_c1_rsr_sft1rstf),
      .cur_rcc_c1_rsr_porrstf  (cur_rcc_c1_rsr_porrstf),
      .cur_rcc_c1_rsr_pinrstf  (cur_rcc_c1_rsr_pinrstf),
      .cur_rcc_c1_rsr_borrstf  (cur_rcc_c1_rsr_borrstf),
      .cur_rcc_c1_rsr_d2rstf   (cur_rcc_c1_rsr_d2rstf),
      .cur_rcc_c1_rsr_d1rstf   (cur_rcc_c1_rsr_d1rstf),
      .cur_rcc_c1_rsr_oblrstf  (cur_rcc_c1_rsr_oblrstf),
      .cur_rcc_c1_rsr_rmvf     (cur_rcc_c1_rsr_rmvf),
      .cur_rcc_c2_rsr_lpwr2rstf(cur_rcc_c2_rsr_lpwr2rstf),
      .cur_rcc_c2_rsr_lpwr1rstf(cur_rcc_c2_rsr_lpwr1rstf),
      .cur_rcc_c2_rsr_wwdg2rstf(cur_rcc_c2_rsr_wwdg2rstf),
      .cur_rcc_c2_rsr_wwdg1rstf(cur_rcc_c2_rsr_wwdg1rstf),
      .cur_rcc_c2_rsr_iwdg2rstf(cur_rcc_c2_rsr_iwdg2rstf),
      .cur_rcc_c2_rsr_iwdg1rstf(cur_rcc_c2_rsr_iwdg1rstf),
      .cur_rcc_c2_rsr_sft2rstf (cur_rcc_c2_rsr_sft2rstf),
      .cur_rcc_c2_rsr_sft1rstf (cur_rcc_c2_rsr_sft1rstf),
      .cur_rcc_c2_rsr_porrstf  (cur_rcc_c2_rsr_porrstf),
      .cur_rcc_c2_rsr_pinrstf  (cur_rcc_c2_rsr_pinrstf),
      .cur_rcc_c2_rsr_borrstf  (cur_rcc_c2_rsr_borrstf),
      .cur_rcc_c2_rsr_d2rstf   (cur_rcc_c2_rsr_d2rstf),
      .cur_rcc_c2_rsr_d1rstf   (cur_rcc_c2_rsr_d1rstf),
      .cur_rcc_c2_rsr_oblrstf  (cur_rcc_c2_rsr_oblrstf),
      .cur_rcc_c2_rsr_rmvf     (cur_rcc_c2_rsr_rmvf),
      .cur_rcc_csr_lsirdy      (cur_rcc_csr_lsirdy),
      .cur_rcc_csr_lsion       (cur_rcc_csr_lsion)
  );

  rcc_vcore_top #(
      .CLK_ON_AFTER_PER_RST_RELEASE (CLK_ON_AFTER_PER_RST_RELEASE),
      .CLK_ON_AFTER_SYS_RST_RELEASE (CLK_ON_AFTER_SYS_RST_RELEASE),
      .CLK_ON_AFTER_D1_RST_RELEASE  (CLK_ON_AFTER_D1_RST_RELEASE),
      .CLK_ON_AFTER_D2_RST_RELEASE  (CLK_ON_AFTER_D2_RST_RELEASE),
      .CLK_ON_AFTER_CPU1_RST_RELEASE(CLK_ON_AFTER_CPU1_RST_RELEASE),
      .CLK_ON_AFTER_CPU2_RST_RELEASE(CLK_ON_AFTER_CPU2_RST_RELEASE)
  ) u_rcc_vcore_top (
      .nrst_in                 (nrst_in),
      .iwdg1_out_rst           (iwdg1_out_rst),
      .wwdg1_out_rst           (wwdg1_out_rst),
      .iwdg2_out_rst           (iwdg2_out_rst),
      .wwdg2_out_rst           (wwdg2_out_rst),
      .lpwr2_rst               (lpwr2_rst),
      .lpwr1_rst               (lpwr1_rst),
      .pwr_bor_rst             (pwr_bor_rst),
      .pwr_por_rst             (pwr_por_rst),
      .cpu2_sftrst             (cpu2_sftrst),
      .cpu1_sftrst             (cpu1_sftrst),
      .d3_deepsleep            (d3_deepsleep),
      .pwr_d1_wkup             (pwr_d1_wkup),
      .pwr_d2_wkup             (pwr_d2_wkup),
      .pwr_d3_wkup             (pwr_d3_wkup),
      .flash_power_ok          (flash_power_ok),
      .pwr_d1_ok               (pwr_d1_ok),
      .pwr_d2_ok               (pwr_d2_ok),
      .pwr_vcore_ok            (pwr_vcore_ok),
      .backup_protect          (backup_protect),
      .c2_sleep                (c2_sleep),
      .c2_deepsleep            (c2_deepsleep),
      .c1_sleep                (c1_sleep),
      .c1_deepsleep            (c1_deepsleep),
      .pad_rcc_eth_mii_tx_clk  (pad_rcc_eth_mii_tx_clk),
      .pad_rcc_eth_mii_rx_clk  (pad_rcc_eth_mii_rx_clk),
      .USB_PHY1                (USB_PHY1),
      .flash_obl_reload        (flash_obl_reload),
      .obl_done                (obl_done),
      .rcc_arcg_on             (rcc_arcg_on),
      .pll3_rdy                (pll3_rdy),
      .pll2_rdy                (pll2_rdy),
      .pll1_rdy                (pll1_rdy),
      .hse_rdy                 (hse_rdy),
      .hsi48_rdy               (hsi48_rdy),
      .csi_rdy                 (csi_rdy),
      .hsi_rdy                 (hsi_rdy),
      .flash_csi_opt           (flash_csi_opt),
      .flash_hsi_opt           (flash_hsi_opt),
      .crs_hsi48_trim          (crs_hsi48_trim),
      .rcc_hsecss_fail         (rcc_hsecss_fail),
      .rcc_lsecss_fail         (rcc_lsecss_fail),
      .ahb_hclk                (ahb_hclk),
      .ahb_hresetn             (ahb_hresetn),
      .ahb_haddr               (ahb_haddr),
      .ahb_hburst              (ahb_hburst),
      .ahb_hprot               (ahb_hprot),
      .ahb_hready_in           (ahb_hready_in),
      .ahb_hsize               (ahb_hsize),
      .ahb_htrans              (ahb_htrans),
      .ahb_hwdata              (ahb_hwdata),
      .ahb_hwrite              (ahb_hwrite),
      .ahb_hsel                (ahb_hsel),
      .ahb_hmaster             (ahb_hmaster),
      .uart8_ker_clk_req       (uart8_ker_clk_req),
      .uart7_ker_clk_req       (uart7_ker_clk_req),
      .i2c3_ker_clk_req        (i2c3_ker_clk_req),
      .i2c2_ker_clk_req        (i2c2_ker_clk_req),
      .i2c1_ker_clk_req        (i2c1_ker_clk_req),
      .uart5_ker_clk_req       (uart5_ker_clk_req),
      .uart4_ker_clk_req       (uart4_ker_clk_req),
      .usart3_ker_clk_req      (usart3_ker_clk_req),
      .usart2_ker_clk_req      (usart2_ker_clk_req),
      .usart6_ker_clk_req      (usart6_ker_clk_req),
      .usart1_ker_clk_req      (usart1_ker_clk_req),
      .i2c4_ker_clk_req        (i2c4_ker_clk_req),
      .lpuart1_ker_clk_req     (lpuart1_ker_clk_req),
      .pll1_p_clk              (pll1_p_clk),
      .pll1_q_clk              (pll1_q_clk),
      .pll2_p_clk              (pll2_p_clk),
      .pll2_q_clk              (pll2_q_clk),
      .pll2_r_clk              (pll2_r_clk),
      .pll3_p_clk              (pll3_p_clk),
      .pll3_q_clk              (pll3_q_clk),
      .pll3_r_clk              (pll3_r_clk),
      .I2S_clk_IN              (I2S_clk_IN),
      .axibridge_d1_busy       (axibridge_d1_busy),
      .ahb3bridge_d1_busy      (ahb3bridge_d1_busy),
      .apb3bridge_d1_busy      (apb3bridge_d1_busy),
      .ahb1bridge_d2_busy      (ahb1bridge_d2_busy),
      .ahb2bridge_d2_busy      (ahb2bridge_d2_busy),
      .apb1bridge_d2_busy      (apb1bridge_d2_busy),
      .apb2bridge_d2_busy      (apb2bridge_d2_busy),
      .ahb4bridge_d3_busy      (ahb4bridge_d3_busy),
      .apb4bridge_d3_busy      (apb4bridge_d3_busy),
      .flash_busy              (flash_busy),
      .hse_css_fail            (hse_css_fail),
      .hse_clk_pre             (hse_clk_pre),
      .lse_clk                 (lse_clk),
      .lsi_clk                 (lsi_clk),
      .hsi48_clk               (hsi48_clk),
      .csi_clk_pre             (csi_clk_pre),
      .hsi_origin_clk          (hsi_origin_clk),
      .eth_rcc_fes             (eth_rcc_fes),
      .eth_rcc_epis_2          (eth_rcc_epis_2),
      .cur_rcc_bdcr_bdrst      (cur_rcc_bdcr_bdrst),
      .cur_rcc_bdcr_rtcen      (cur_rcc_bdcr_rtcen),
      .cur_rcc_bdcr_rtcsel     (cur_rcc_bdcr_rtcsel),
      .cur_rcc_bdcr_lsecssd    (cur_rcc_bdcr_lsecssd),
      .cur_rcc_bdcr_lsecsson   (cur_rcc_bdcr_lsecsson),
      .cur_rcc_bdcr_lsedrv     (cur_rcc_bdcr_lsedrv),
      .cur_rcc_bdcr_lsebyp     (cur_rcc_bdcr_lsebyp),
      .cur_rcc_bdcr_lserdy     (cur_rcc_bdcr_lserdy),
      .cur_rcc_bdcr_lseon      (cur_rcc_bdcr_lseon),
      .cur_rcc_c1_rsr_lpwr2rstf(cur_rcc_c1_rsr_lpwr2rstf),
      .cur_rcc_c1_rsr_lpwr1rstf(cur_rcc_c1_rsr_lpwr1rstf),
      .cur_rcc_c1_rsr_wwdg2rstf(cur_rcc_c1_rsr_wwdg2rstf),
      .cur_rcc_c1_rsr_wwdg1rstf(cur_rcc_c1_rsr_wwdg1rstf),
      .cur_rcc_c1_rsr_iwdg2rstf(cur_rcc_c1_rsr_iwdg2rstf),
      .cur_rcc_c1_rsr_iwdg1rstf(cur_rcc_c1_rsr_iwdg1rstf),
      .cur_rcc_c1_rsr_sft2rstf (cur_rcc_c1_rsr_sft2rstf),
      .cur_rcc_c1_rsr_sft1rstf (cur_rcc_c1_rsr_sft1rstf),
      .cur_rcc_c1_rsr_porrstf  (cur_rcc_c1_rsr_porrstf),
      .cur_rcc_c1_rsr_pinrstf  (cur_rcc_c1_rsr_pinrstf),
      .cur_rcc_c1_rsr_borrstf  (cur_rcc_c1_rsr_borrstf),
      .cur_rcc_c1_rsr_d2rstf   (cur_rcc_c1_rsr_d2rstf),
      .cur_rcc_c1_rsr_d1rstf   (cur_rcc_c1_rsr_d1rstf),
      .cur_rcc_c1_rsr_oblrstf  (cur_rcc_c1_rsr_oblrstf),
      .cur_rcc_c1_rsr_rmvf     (cur_rcc_c1_rsr_rmvf),
      .cur_rcc_c2_rsr_lpwr2rstf(cur_rcc_c2_rsr_lpwr2rstf),
      .cur_rcc_c2_rsr_lpwr1rstf(cur_rcc_c2_rsr_lpwr1rstf),
      .cur_rcc_c2_rsr_wwdg2rstf(cur_rcc_c2_rsr_wwdg2rstf),
      .cur_rcc_c2_rsr_wwdg1rstf(cur_rcc_c2_rsr_wwdg1rstf),
      .cur_rcc_c2_rsr_iwdg2rstf(cur_rcc_c2_rsr_iwdg2rstf),
      .cur_rcc_c2_rsr_iwdg1rstf(cur_rcc_c2_rsr_iwdg1rstf),
      .cur_rcc_c2_rsr_sft2rstf (cur_rcc_c2_rsr_sft2rstf),
      .cur_rcc_c2_rsr_sft1rstf (cur_rcc_c2_rsr_sft1rstf),
      .cur_rcc_c2_rsr_porrstf  (cur_rcc_c2_rsr_porrstf),
      .cur_rcc_c2_rsr_pinrstf  (cur_rcc_c2_rsr_pinrstf),
      .cur_rcc_c2_rsr_borrstf  (cur_rcc_c2_rsr_borrstf),
      .cur_rcc_c2_rsr_d2rstf   (cur_rcc_c2_rsr_d2rstf),
      .cur_rcc_c2_rsr_d1rstf   (cur_rcc_c2_rsr_d1rstf),
      .cur_rcc_c2_rsr_oblrstf  (cur_rcc_c2_rsr_oblrstf),
      .cur_rcc_c2_rsr_rmvf     (cur_rcc_c2_rsr_rmvf),
      .cur_rcc_csr_lsirdy      (cur_rcc_csr_lsirdy),
      .cur_rcc_csr_lsion       (cur_rcc_csr_lsion),

      .nrst_out                 (nrst_out),
      .rcc_pwr_d1_req           (rcc_pwr_d1_req),
      .rcc_pwr_d2_req           (rcc_pwr_d2_req),
      .rcc_pwr_d3_req           (rcc_pwr_d3_req),
      .c2_per_alloc_d1          (c2_per_alloc_d1),
      .c1_per_alloc_d2          (c1_per_alloc_d2),
      .rcc_c2_clk               (rcc_c2_clk),
      .rcc_fclk_c2              (rcc_fclk_c2),
      .rcc_c2_systick_clk       (rcc_c2_systick_clk),
      .rcc_c1_clk               (rcc_c1_clk),
      .rcc_fclk_c1              (rcc_fclk_c1),
      .rcc_c1_systick_clk       (rcc_c1_systick_clk),
      .cpu1_arcg_rst_n          (cpu1_arcg_rst_n),
      .cpu2_arcg_rst_n          (cpu2_arcg_rst_n),
      .d1_bus_arcg_rst_n        (d1_bus_arcg_rst_n),
      .d2_bus_arcg_rst_n        (d2_bus_arcg_rst_n),
      .d3_bus_arcg_rst_n        (d3_bus_arcg_rst_n),
      .rcc_timx_ker_clk         (rcc_timx_ker_clk),
      .rcc_timy_ker_clk         (rcc_timy_ker_clk),
      .rcc_hrtimer_prescalar_clk(rcc_hrtimer_prescalar_clk),
      .sys_d1cpre_clk           (sys_d1cpre_clk),
      .sys_hpre_clk             (sys_hpre_clk),
      .hse_rtc_clk              (hse_rtc_clk),
      .mco1                     (mco1),
      .mco2                     (mco2),
      .rcc_hsefail_it           (rcc_hsefail_it),
      .rcc_lsefail_it           (rcc_lsefail_it),
      .rcc_it                   (rcc_it),
      .pwr_por_rst_n            (pwr_por_rst_n),
      .sys_arcg_rst_n           (sys_arcg_rst_n),
      .d1_arcg_rst_n            (d1_arcg_rst_n),
      .d2_arcg_rst_n            (d2_arcg_rst_n),
      .stby_rst_n               (stby_rst_n),
      .rcc_flash_arcg_rst_n     (rcc_flash_arcg_rst_n),
      .rcc_qspi_arcg_rst_n      (rcc_qspi_arcg_rst_n),
      .rcc_axisram_arcg_rst_n   (rcc_axisram_arcg_rst_n),
      .rcc_fmc_arcg_rst_n       (rcc_fmc_arcg_rst_n),
      .rcc_dma2d_arcg_rst_n     (rcc_dma2d_arcg_rst_n),
      .rcc_mdma_arcg_rst_n      (rcc_mdma_arcg_rst_n),
      .rcc_ltdc_arcg_rst_n      (rcc_ltdc_arcg_rst_n),
      .rcc_ramecc1_arcg_rst_n   (rcc_ramecc1_arcg_rst_n),
      .rcc_gpv_arcg_rst_n       (rcc_gpv_arcg_rst_n),
      .rcc_itcm_arcg_rst_n      (rcc_itcm_arcg_rst_n),
      .rcc_dtcm2_arcg_rst_n     (rcc_dtcm2_arcg_rst_n),
      .rcc_dtcm1_arcg_rst_n     (rcc_dtcm1_arcg_rst_n),
      .rcc_jpgdec_arcg_rst_n    (rcc_jpgdec_arcg_rst_n),
      .rcc_sdmmc1_arcg_rst_n    (rcc_sdmmc1_arcg_rst_n),
      .rcc_wwdg1_arcg_rst_n     (rcc_wwdg1_arcg_rst_n),
      .rcc_usb2ulpi_arcg_rst_n  (rcc_usb2ulpi_arcg_rst_n),
      .rcc_usb2otg_arcg_rst_n   (rcc_usb2otg_arcg_rst_n),
      .rcc_usb1ulpi_arcg_rst_n  (rcc_usb1ulpi_arcg_rst_n),
      .rcc_usb1otg_arcg_rst_n   (rcc_usb1otg_arcg_rst_n),
      .rcc_eth1rx_arcg_rst_n    (rcc_eth1rx_arcg_rst_n),
      .rcc_eth1tx_arcg_rst_n    (rcc_eth1tx_arcg_rst_n),
      .rcc_eth1mac_arcg_rst_n   (rcc_eth1mac_arcg_rst_n),
      .rcc_adc12_arcg_rst_n     (rcc_adc12_arcg_rst_n),
      .rcc_dma2_arcg_rst_n      (rcc_dma2_arcg_rst_n),
      .rcc_dma1_arcg_rst_n      (rcc_dma1_arcg_rst_n),
      .rcc_sram3_arcg_rst_n     (rcc_sram3_arcg_rst_n),
      .rcc_sram2_arcg_rst_n     (rcc_sram2_arcg_rst_n),
      .rcc_sram1_arcg_rst_n     (rcc_sram1_arcg_rst_n),
      .rcc_sdmmc2_arcg_rst_n    (rcc_sdmmc2_arcg_rst_n),
      .rcc_rng_arcg_rst_n       (rcc_rng_arcg_rst_n),
      .rcc_hash_arcg_rst_n      (rcc_hash_arcg_rst_n),
      .rcc_crypt_arcg_rst_n     (rcc_crypt_arcg_rst_n),
      .rcc_dcmi_arcg_rst_n      (rcc_dcmi_arcg_rst_n),
      .rcc_ramecc2_arcg_rst_n   (rcc_ramecc2_arcg_rst_n),
      .rcc_uart8_arcg_rst_n     (rcc_uart8_arcg_rst_n),
      .rcc_uart7_arcg_rst_n     (rcc_uart7_arcg_rst_n),
      .rcc_dac12_arcg_rst_n     (rcc_dac12_arcg_rst_n),
      .rcc_hdmicec_arcg_rst_n   (rcc_hdmicec_arcg_rst_n),
      .rcc_i2c3_arcg_rst_n      (rcc_i2c3_arcg_rst_n),
      .rcc_i2c2_arcg_rst_n      (rcc_i2c2_arcg_rst_n),
      .rcc_i2c1_arcg_rst_n      (rcc_i2c1_arcg_rst_n),
      .rcc_uart5_arcg_rst_n     (rcc_uart5_arcg_rst_n),
      .rcc_uart4_arcg_rst_n     (rcc_uart4_arcg_rst_n),
      .rcc_usart3_arcg_rst_n    (rcc_usart3_arcg_rst_n),
      .rcc_usart2_arcg_rst_n    (rcc_usart2_arcg_rst_n),
      .rcc_spdifrx_arcg_rst_n   (rcc_spdifrx_arcg_rst_n),
      .rcc_spi3_arcg_rst_n      (rcc_spi3_arcg_rst_n),
      .rcc_spi2_arcg_rst_n      (rcc_spi2_arcg_rst_n),
      .rcc_wwdg2_arcg_rst_n     (rcc_wwdg2_arcg_rst_n),
      .rcc_lptim1_arcg_rst_n    (rcc_lptim1_arcg_rst_n),
      .rcc_tim14_arcg_rst_n     (rcc_tim14_arcg_rst_n),
      .rcc_tim13_arcg_rst_n     (rcc_tim13_arcg_rst_n),
      .rcc_tim12_arcg_rst_n     (rcc_tim12_arcg_rst_n),
      .rcc_tim7_arcg_rst_n      (rcc_tim7_arcg_rst_n),
      .rcc_tim6_arcg_rst_n      (rcc_tim6_arcg_rst_n),
      .rcc_tim5_arcg_rst_n      (rcc_tim5_arcg_rst_n),
      .rcc_tim4_arcg_rst_n      (rcc_tim4_arcg_rst_n),
      .rcc_tim3_arcg_rst_n      (rcc_tim3_arcg_rst_n),
      .rcc_tim2_arcg_rst_n      (rcc_tim2_arcg_rst_n),
      .rcc_fdcan_arcg_rst_n     (rcc_fdcan_arcg_rst_n),
      .rcc_mdios_arcg_rst_n     (rcc_mdios_arcg_rst_n),
      .rcc_opamp_arcg_rst_n     (rcc_opamp_arcg_rst_n),
      .rcc_swpmi_arcg_rst_n     (rcc_swpmi_arcg_rst_n),
      .rcc_crs_arcg_rst_n       (rcc_crs_arcg_rst_n),
      .rcc_hrtim_arcg_rst_n     (rcc_hrtim_arcg_rst_n),
      .rcc_dfsdm1_arcg_rst_n    (rcc_dfsdm1_arcg_rst_n),
      .rcc_sai3_arcg_rst_n      (rcc_sai3_arcg_rst_n),
      .rcc_sai2_arcg_rst_n      (rcc_sai2_arcg_rst_n),
      .rcc_sai1_arcg_rst_n      (rcc_sai1_arcg_rst_n),
      .rcc_spi5_arcg_rst_n      (rcc_spi5_arcg_rst_n),
      .rcc_tim17_arcg_rst_n     (rcc_tim17_arcg_rst_n),
      .rcc_tim16_arcg_rst_n     (rcc_tim16_arcg_rst_n),
      .rcc_tim15_arcg_rst_n     (rcc_tim15_arcg_rst_n),
      .rcc_spi4_arcg_rst_n      (rcc_spi4_arcg_rst_n),
      .rcc_spi1_arcg_rst_n      (rcc_spi1_arcg_rst_n),
      .rcc_usart6_arcg_rst_n    (rcc_usart6_arcg_rst_n),
      .rcc_usart1_arcg_rst_n    (rcc_usart1_arcg_rst_n),
      .rcc_tim8_arcg_rst_n      (rcc_tim8_arcg_rst_n),
      .rcc_tim1_arcg_rst_n      (rcc_tim1_arcg_rst_n),
      .rcc_sram4_arcg_rst_n     (rcc_sram4_arcg_rst_n),
      .rcc_bkpram_arcg_rst_n    (rcc_bkpram_arcg_rst_n),
      .rcc_ramecc3_arcg_rst_n   (rcc_ramecc3_arcg_rst_n),
      .rcc_hsem_arcg_rst_n      (rcc_hsem_arcg_rst_n),
      .rcc_adc3_arcg_rst_n      (rcc_adc3_arcg_rst_n),
      .rcc_bdma_arcg_rst_n      (rcc_bdma_arcg_rst_n),
      .rcc_crc_arcg_rst_n       (rcc_crc_arcg_rst_n),
      .rcc_gpiok_arcg_rst_n     (rcc_gpiok_arcg_rst_n),
      .rcc_gpioj_arcg_rst_n     (rcc_gpioj_arcg_rst_n),
      .rcc_gpioi_arcg_rst_n     (rcc_gpioi_arcg_rst_n),
      .rcc_gpioh_arcg_rst_n     (rcc_gpioh_arcg_rst_n),
      .rcc_gpiog_arcg_rst_n     (rcc_gpiog_arcg_rst_n),
      .rcc_gpiof_arcg_rst_n     (rcc_gpiof_arcg_rst_n),
      .rcc_gpioe_arcg_rst_n     (rcc_gpioe_arcg_rst_n),
      .rcc_gpiod_arcg_rst_n     (rcc_gpiod_arcg_rst_n),
      .rcc_gpioc_arcg_rst_n     (rcc_gpioc_arcg_rst_n),
      .rcc_gpiob_arcg_rst_n     (rcc_gpiob_arcg_rst_n),
      .rcc_gpioa_arcg_rst_n     (rcc_gpioa_arcg_rst_n),
      .rcc_rcc_arcg_rst_n       (rcc_rcc_arcg_rst_n),
      .rcc_pwr_arcg_rst_n       (rcc_pwr_arcg_rst_n),
      .rcc_sai4_arcg_rst_n      (rcc_sai4_arcg_rst_n),
      .rcc_rtc_arcg_rst_n       (rcc_rtc_arcg_rst_n),
      .rcc_vref_arcg_rst_n      (rcc_vref_arcg_rst_n),
      .rcc_comp12_arcg_rst_n    (rcc_comp12_arcg_rst_n),
      .rcc_lptim5_arcg_rst_n    (rcc_lptim5_arcg_rst_n),
      .rcc_lptim4_arcg_rst_n    (rcc_lptim4_arcg_rst_n),
      .rcc_lptim3_arcg_rst_n    (rcc_lptim3_arcg_rst_n),
      .rcc_lptim2_arcg_rst_n    (rcc_lptim2_arcg_rst_n),
      .rcc_i2c4_arcg_rst_n      (rcc_i2c4_arcg_rst_n),
      .rcc_spi6_arcg_rst_n      (rcc_spi6_arcg_rst_n),
      .rcc_lpuart1_arcg_rst_n   (rcc_lpuart1_arcg_rst_n),
      .rcc_syscfg_arcg_rst_n    (rcc_syscfg_arcg_rst_n),
      .rcc_iwdg2_arcg_rst_n     (rcc_iwdg2_arcg_rst_n),
      .rcc_iwdg1_arcg_rst_n     (rcc_iwdg1_arcg_rst_n),
      .rcc_exti_arcg_rst_n      (rcc_exti_arcg_rst_n),
      .ahb_hrdata               (ahb_hrdata),
      .ahb_hready_out           (ahb_hready_out),
      .ahb_hresp                (ahb_hresp),
      .rcc_axibridge_d1_clk     (rcc_axibridge_d1_clk),
      .rcc_ahb3bridge_d1_clk    (rcc_ahb3bridge_d1_clk),
      .rcc_apb3bridge_d1_clk    (rcc_apb3bridge_d1_clk),
      .rcc_ahb1bridge_d2_clk    (rcc_ahb1bridge_d2_clk),
      .rcc_ahb2bridge_d2_clk    (rcc_ahb2bridge_d2_clk),
      .rcc_apb1bridge_d2_clk    (rcc_apb1bridge_d2_clk),
      .rcc_apb2bridge_d2_clk    (rcc_apb2bridge_d2_clk),
      .rcc_ahb4bridge_d3_clk    (rcc_ahb4bridge_d3_clk),
      .rcc_apb4bridge_d3_clk    (rcc_apb4bridge_d3_clk),
      .pll1_src_clk             (pll1_src_clk),
      .pll2_src_clk             (pll2_src_clk),
      .pll3_src_clk             (pll3_src_clk),
      .pll3on                   (pll3on),
      .pll2on                   (pll2on),
      .pll1on                   (pll1on),
      .hsecsson                 (hsecsson),
      .hsebyp                   (hsebyp),
      .hseon                    (hseon),
      .hsi48on                  (hsi48on),
      .csikeron                 (csikeron),
      .csion                    (csion),
      .hsidiv                   (hsidiv),
      .hsikeron                 (hsikeron),
      .hsion                    (hsion),
      .rcc_csi_triming          (rcc_csi_triming),
      .rcc_hsi_triming          (rcc_hsi_triming),
      .divr3en                  (divr3en),
      .divq3en                  (divq3en),
      .divp3en                  (divp3en),
      .divr2en                  (divr2en),
      .divq2en                  (divq2en),
      .divp2en                  (divp2en),
      .divr1en                  (divr1en),
      .divq1en                  (divq1en),
      .divp1en                  (divp1en),
      .pll3rge                  (pll3rge),
      .pll3vcosel               (pll3vcosel),
      .pll3fracen               (pll3fracen),
      .pll2rge                  (pll2rge),
      .pll2vcosel               (pll2vcosel),
      .pll2fracen               (pll2fracen),
      .pll1rge                  (pll1rge),
      .pll1vcosel               (pll1vcosel),
      .pll1fracen               (pll1fracen),
      .divr1                    (divr1),
      .divq1                    (divq1),
      .divp1                    (divp1),
      .divn1                    (divn1),
      .fracn1                   (fracn1),
      .divr2                    (divr2),
      .divq2                    (divq2),
      .divp2                    (divp2),
      .divn2                    (divn2),
      .fracn2                   (fracn2),
      .divr3                    (divr3),
      .divq3                    (divq3),
      .divp3                    (divp3),
      .divn3                    (divn3),
      .fracn3                   (fracn3),
      .rcc_eth_mii_tx_clk       (rcc_eth_mii_tx_clk),
      .rcc_eth_mii_rx_clk       (rcc_eth_mii_rx_clk),
      .rcc_eth_rmii_ref_clk     (rcc_eth_rmii_ref_clk),
      .rcc_c1_rsr_rmvf_wren     (rcc_c1_rsr_rmvf_wren),
      .rcc_c2_rsr_rmvf_wren     (rcc_c2_rsr_rmvf_wren),
      .rcc_csr_lsion_wren       (rcc_csr_lsion_wren),
      .rcc_bdcr_byte2_wren      (rcc_bdcr_byte2_wren),
      .rcc_bdcr_byte1_wren      (rcc_bdcr_byte1_wren),
      .rcc_bdcr_byte0_wren      (rcc_bdcr_byte0_wren),
      .nxt_rcc_bdcr_bdrst       (nxt_rcc_bdcr_bdrst),
      .nxt_rcc_bdcr_rtcen       (nxt_rcc_bdcr_rtcen),
      .nxt_rcc_bdcr_rtcsel      (nxt_rcc_bdcr_rtcsel),
      .nxt_rcc_bdcr_lsecsson    (nxt_rcc_bdcr_lsecsson),
      .nxt_rcc_bdcr_lsedrv      (nxt_rcc_bdcr_lsedrv),
      .nxt_rcc_bdcr_lsebyp      (nxt_rcc_bdcr_lsebyp),
      .nxt_rcc_bdcr_lseon       (nxt_rcc_bdcr_lseon),
      .rcc_rtc_pclk             (rcc_rtc_pclk),
      .rcc_flash_aclk           (rcc_flash_aclk),
      .rcc_flash_hclk           (rcc_flash_hclk),
      .rcc_qspi_aclk            (rcc_qspi_aclk),
      .rcc_qspi_hclk            (rcc_qspi_hclk),
      .rcc_qspi_ker_clk         (rcc_qspi_ker_clk),
      .rcc_axisram_aclk         (rcc_axisram_aclk),
      .rcc_fmc_aclk             (rcc_fmc_aclk),
      .rcc_fmc_hclk             (rcc_fmc_hclk),
      .rcc_fmc_ker_clk          (rcc_fmc_ker_clk),
      .rcc_dma2d_aclk           (rcc_dma2d_aclk),
      .rcc_dma2d_hclk           (rcc_dma2d_hclk),
      .rcc_mdma_aclk            (rcc_mdma_aclk),
      .rcc_mdma_hclk            (rcc_mdma_hclk),
      .rcc_ltdc_aclk            (rcc_ltdc_aclk),
      .rcc_ltdc_pclk            (rcc_ltdc_pclk),
      .rcc_ltdc_ker_clk         (rcc_ltdc_ker_clk),
      .rcc_ramecc1_hclk         (rcc_ramecc1_hclk),
      .rcc_gpv_hclk             (rcc_gpv_hclk),
      .rcc_itcm_hclk            (rcc_itcm_hclk),
      .rcc_dtcm2_hclk           (rcc_dtcm2_hclk),
      .rcc_dtcm1_hclk           (rcc_dtcm1_hclk),
      .rcc_jpgdec_hclk          (rcc_jpgdec_hclk),
      .rcc_sdmmc1_hclk          (rcc_sdmmc1_hclk),
      .rcc_sdmmc1_ker_clk       (rcc_sdmmc1_ker_clk),
      .rcc_wwdg1_pclk           (rcc_wwdg1_pclk),
      .rcc_usb2ulpi_hclk        (rcc_usb2ulpi_hclk),
      .rcc_usb2otg_hclk         (rcc_usb2otg_hclk),
      .rcc_usb2otg_ker_clk      (rcc_usb2otg_ker_clk),
      .rcc_usb1ulpi_hclk        (rcc_usb1ulpi_hclk),
      .rcc_usb1ulpi_ker_clk     (rcc_usb1ulpi_ker_clk),
      .rcc_usb1otg_hclk         (rcc_usb1otg_hclk),
      .rcc_usb1otg_ker_clk      (rcc_usb1otg_ker_clk),
      .rcc_eth1rx_hclk          (rcc_eth1rx_hclk),
      .rcc_eth1tx_hclk          (rcc_eth1tx_hclk),
      .rcc_eth1mac_hclk         (rcc_eth1mac_hclk),
      .rcc_adc12_hclk           (rcc_adc12_hclk),
      .rcc_adc12_ker_clk        (rcc_adc12_ker_clk),
      .rcc_dma2_hclk            (rcc_dma2_hclk),
      .rcc_dma1_hclk            (rcc_dma1_hclk),
      .rcc_sram3_hclk           (rcc_sram3_hclk),
      .rcc_sram2_hclk           (rcc_sram2_hclk),
      .rcc_sram1_hclk           (rcc_sram1_hclk),
      .rcc_sdmmc2_hclk          (rcc_sdmmc2_hclk),
      .rcc_sdmmc2_ker_clk       (rcc_sdmmc2_ker_clk),
      .rcc_rng_hclk             (rcc_rng_hclk),
      .rcc_rng_ker_clk          (rcc_rng_ker_clk),
      .rcc_hash_hclk            (rcc_hash_hclk),
      .rcc_crypt_hclk           (rcc_crypt_hclk),
      .rcc_dcmi_hclk            (rcc_dcmi_hclk),
      .rcc_ramecc2_hclk         (rcc_ramecc2_hclk),
      .rcc_uart8_pclk           (rcc_uart8_pclk),
      .rcc_uart8_ker_clk        (rcc_uart8_ker_clk),
      .rcc_uart7_pclk           (rcc_uart7_pclk),
      .rcc_uart7_ker_clk        (rcc_uart7_ker_clk),
      .rcc_dac12_pclk           (rcc_dac12_pclk),
      .rcc_hdmicec_pclk         (rcc_hdmicec_pclk),
      .rcc_hdmicec_ker_clk      (rcc_hdmicec_ker_clk),
      .rcc_i2c3_pclk            (rcc_i2c3_pclk),
      .rcc_i2c3_ker_clk         (rcc_i2c3_ker_clk),
      .rcc_i2c2_pclk            (rcc_i2c2_pclk),
      .rcc_i2c2_ker_clk         (rcc_i2c2_ker_clk),
      .rcc_i2c1_pclk            (rcc_i2c1_pclk),
      .rcc_i2c1_ker_clk         (rcc_i2c1_ker_clk),
      .rcc_uart5_pclk           (rcc_uart5_pclk),
      .rcc_uart5_ker_clk        (rcc_uart5_ker_clk),
      .rcc_uart4_pclk           (rcc_uart4_pclk),
      .rcc_uart4_ker_clk        (rcc_uart4_ker_clk),
      .rcc_usart3_pclk          (rcc_usart3_pclk),
      .rcc_usart3_ker_clk       (rcc_usart3_ker_clk),
      .rcc_usart2_pclk          (rcc_usart2_pclk),
      .rcc_usart2_ker_clk       (rcc_usart2_ker_clk),
      .rcc_spdifrx_pclk         (rcc_spdifrx_pclk),
      .rcc_spdifrx_ker_clk      (rcc_spdifrx_ker_clk),
      .rcc_spi3_pclk            (rcc_spi3_pclk),
      .rcc_spi3_ker_clk         (rcc_spi3_ker_clk),
      .rcc_spi2_pclk            (rcc_spi2_pclk),
      .rcc_spi2_ker_clk         (rcc_spi2_ker_clk),
      .rcc_wwdg2_pclk           (rcc_wwdg2_pclk),
      .rcc_lptim1_pclk          (rcc_lptim1_pclk),
      .rcc_lptim1_ker_clk       (rcc_lptim1_ker_clk),
      .rcc_tim14_pclk           (rcc_tim14_pclk),
      .rcc_tim14_ker_clk        (rcc_tim14_ker_clk),
      .rcc_tim13_pclk           (rcc_tim13_pclk),
      .rcc_tim13_ker_clk        (rcc_tim13_ker_clk),
      .rcc_tim12_pclk           (rcc_tim12_pclk),
      .rcc_tim12_ker_clk        (rcc_tim12_ker_clk),
      .rcc_tim7_pclk            (rcc_tim7_pclk),
      .rcc_tim7_ker_clk         (rcc_tim7_ker_clk),
      .rcc_tim6_pclk            (rcc_tim6_pclk),
      .rcc_tim6_ker_clk         (rcc_tim6_ker_clk),
      .rcc_tim5_pclk            (rcc_tim5_pclk),
      .rcc_tim5_ker_clk         (rcc_tim5_ker_clk),
      .rcc_tim4_pclk            (rcc_tim4_pclk),
      .rcc_tim4_ker_clk         (rcc_tim4_ker_clk),
      .rcc_tim3_pclk            (rcc_tim3_pclk),
      .rcc_tim3_ker_clk         (rcc_tim3_ker_clk),
      .rcc_tim2_pclk            (rcc_tim2_pclk),
      .rcc_tim2_ker_clk         (rcc_tim2_ker_clk),
      .rcc_fdcan_pclk           (rcc_fdcan_pclk),
      .rcc_fdcan_ker_clk        (rcc_fdcan_ker_clk),
      .rcc_mdios_pclk           (rcc_mdios_pclk),
      .rcc_opamp_pclk           (rcc_opamp_pclk),
      .rcc_swpmi_pclk           (rcc_swpmi_pclk),
      .rcc_swpmi_ker_clk        (rcc_swpmi_ker_clk),
      .rcc_crs_pclk             (rcc_crs_pclk),
      .rcc_hrtim_pclk           (rcc_hrtim_pclk),
      .rcc_hrtim_ker_clk        (rcc_hrtim_ker_clk),
      .rcc_dfsdm1_pclk          (rcc_dfsdm1_pclk),
      .rcc_dfsdm1_ker_clk_0     (rcc_dfsdm1_ker_clk_0),
      .rcc_dfsdm1_ker_clk_1     (rcc_dfsdm1_ker_clk_1),
      .rcc_sai3_pclk            (rcc_sai3_pclk),
      .rcc_sai3_ker_clk         (rcc_sai3_ker_clk),
      .rcc_sai2_pclk            (rcc_sai2_pclk),
      .rcc_sai2_ker_clk         (rcc_sai2_ker_clk),
      .rcc_sai1_pclk            (rcc_sai1_pclk),
      .rcc_sai1_ker_clk         (rcc_sai1_ker_clk),
      .rcc_spi5_pclk            (rcc_spi5_pclk),
      .rcc_spi5_ker_clk         (rcc_spi5_ker_clk),
      .rcc_tim17_pclk           (rcc_tim17_pclk),
      .rcc_tim17_ker_clk        (rcc_tim17_ker_clk),
      .rcc_tim16_pclk           (rcc_tim16_pclk),
      .rcc_tim16_ker_clk        (rcc_tim16_ker_clk),
      .rcc_tim15_pclk           (rcc_tim15_pclk),
      .rcc_tim15_ker_clk        (rcc_tim15_ker_clk),
      .rcc_spi4_pclk            (rcc_spi4_pclk),
      .rcc_spi4_ker_clk         (rcc_spi4_ker_clk),
      .rcc_spi1_pclk            (rcc_spi1_pclk),
      .rcc_spi1_ker_clk         (rcc_spi1_ker_clk),
      .rcc_usart6_pclk          (rcc_usart6_pclk),
      .rcc_usart6_ker_clk       (rcc_usart6_ker_clk),
      .rcc_usart1_pclk          (rcc_usart1_pclk),
      .rcc_usart1_ker_clk       (rcc_usart1_ker_clk),
      .rcc_tim8_pclk            (rcc_tim8_pclk),
      .rcc_tim8_ker_clk         (rcc_tim8_ker_clk),
      .rcc_tim1_pclk            (rcc_tim1_pclk),
      .rcc_tim1_ker_clk         (rcc_tim1_ker_clk),
      .rcc_sram4_hclk           (rcc_sram4_hclk),
      .rcc_bkpram_hclk          (rcc_bkpram_hclk),
      .rcc_ramecc3_hclk         (rcc_ramecc3_hclk),
      .rcc_hsem_hclk            (rcc_hsem_hclk),
      .rcc_adc3_hclk            (rcc_adc3_hclk),
      .rcc_adc3_ker_clk         (rcc_adc3_ker_clk),
      .rcc_bdma_hclk            (rcc_bdma_hclk),
      .rcc_crc_hclk             (rcc_crc_hclk),
      .rcc_gpiok_hclk           (rcc_gpiok_hclk),
      .rcc_gpioj_hclk           (rcc_gpioj_hclk),
      .rcc_gpioi_hclk           (rcc_gpioi_hclk),
      .rcc_gpioh_hclk           (rcc_gpioh_hclk),
      .rcc_gpiog_hclk           (rcc_gpiog_hclk),
      .rcc_gpiof_hclk           (rcc_gpiof_hclk),
      .rcc_gpioe_hclk           (rcc_gpioe_hclk),
      .rcc_gpiod_hclk           (rcc_gpiod_hclk),
      .rcc_gpioc_hclk           (rcc_gpioc_hclk),
      .rcc_gpiob_hclk           (rcc_gpiob_hclk),
      .rcc_gpioa_hclk           (rcc_gpioa_hclk),
      .rcc_rcc_hclk             (rcc_rcc_hclk),
      .rcc_pwr_hclk             (rcc_pwr_hclk),
      .rcc_sai4_pclk            (rcc_sai4_pclk),
      .rcc_sai4_ker_clk_0       (rcc_sai4_ker_clk_0),
      .rcc_sai4_ker_clk_1       (rcc_sai4_ker_clk_1),
      .rcc_vref_pclk            (rcc_vref_pclk),
      .rcc_comp12_pclk          (rcc_comp12_pclk),
      .rcc_lptim5_pclk          (rcc_lptim5_pclk),
      .rcc_lptim5_ker_clk       (rcc_lptim5_ker_clk),
      .rcc_lptim4_pclk          (rcc_lptim4_pclk),
      .rcc_lptim4_ker_clk       (rcc_lptim4_ker_clk),
      .rcc_lptim3_pclk          (rcc_lptim3_pclk),
      .rcc_lptim3_ker_clk       (rcc_lptim3_ker_clk),
      .rcc_lptim2_pclk          (rcc_lptim2_pclk),
      .rcc_lptim2_ker_clk       (rcc_lptim2_ker_clk),
      .rcc_i2c4_pclk            (rcc_i2c4_pclk),
      .rcc_i2c4_ker_clk         (rcc_i2c4_ker_clk),
      .rcc_spi6_pclk            (rcc_spi6_pclk),
      .rcc_spi6_ker_clk         (rcc_spi6_ker_clk),
      .rcc_lpuart1_pclk         (rcc_lpuart1_pclk),
      .rcc_lpuart1_ker_clk      (rcc_lpuart1_ker_clk),
      .rcc_syscfg_pclk          (rcc_syscfg_pclk),
      .rcc_iwdg2_pclk           (rcc_iwdg2_pclk),
      .rcc_iwdg1_pclk           (rcc_iwdg1_pclk),
      .rcc_exti_pclk            (rcc_exti_pclk)
  );



endmodule
