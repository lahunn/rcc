module BB_clk_div_d #(
    parameter RATIO_WID = 8
) (
    input  rst_n,
    input  i_clk,
    input  ratio,
    output o_clk,
    output div_en
);
// NULL MODULE

endmodule  //moduleName
