module BB_clk_div_s #(
    parameter DIV_RATIO = 3
) (
    input  rst_n,
    input  i_clk,
    output o_clk,
    output div_en
);
// NULL MODULE


endmodule  //moduleName
