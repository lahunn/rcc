/* verilator lint_off UNUSEDPARAM */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off UNDRIVEN */
module BB_clk_div_s #(
    parameter DIV_RATIO = 3
) (
    input  rst_n,
    input  i_clk,
    output o_clk,
    input  div_en
);
// NULL MODULE


endmodule  //moduleName
