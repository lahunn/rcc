module rcc_top #(
    // parameter D1_AXI_NUM = 1,   // IN NEXT VERSION.we will add these parameter
    // parameter D1_AHB_NUM = 1,
    // parameter D1_APB_NUM = 1,
    // parameter D2_AXI_NUM = 0,
    // parameter D2_AHB_NUM = 2,
    // parameter D2_APB_NUM = 2,
    // parameter D3_AXI_NUM = 0,
    // parameter D3_AHB_NUM = 1,
    // parameter D3_APB_NUM = 1,
    parameter D1_AXI_PER_NUM = 10,
    parameter D1_AHB_PER_NUM = 10,
    parameter D1_APB_PER_NUM = 10,
    parameter D2_AXI_PER_NUM = 0,
    parameter D2_AHB_PER_NUM = 10,
    parameter D2_APB_PER_NUM = 10,
    parameter D3_AXI_PER_NUM = 0,
    parameter D3_AHB_PER_NUM = 10,
    parameter D3_APB_PER_NUM = 10
)( 
// signals connected to PAD 
    input [0:0] OSC32_IN,
    output [0:0] OSC32_OUT,
    input [0:0] OSC_IN,
    output [0:0] OSC_OUT,
    output [0:0] MCO1,
    output [0:0] MCO2,
    input [0:0] ARCG_ON,
    input [0:0] I2S_CLKIN,
    input [0:0] ETH_MII_TX_CLK,
    input [0:0] ETH_MII_RX_CLK,
    input [0:0] ETH_RMII_REF_CLK,
    input [0:0] USB_PHY1,
    input [0:0] USB_PHY2,
// signals connected to PAD_NRST 
    input [0:0] nrst_in,
    output [0:0] nrst_out,
// signals connected to PWR 
    input [0:0] d3_deepsleep,
    input [0:0] pwr_d1_wkup,
    input [0:0] pwr_d2_wkup,
    input [0:0] pwr_d3_wkup,
    output [0:0] rcc_pwd_d1_req,
    output [0:0] rcc_pwd_d2_req,
    output [0:0] rcc_pwd_d3_req,
    output [0:0] cpu_per_alloc_d1,
    output [0:0] cpu_per_alloc_d2,
    input [0:0] flash_power_ok,
    input [0:0] pwr_d1_ok,
    input [0:0] pwr_d2_ok,
    input [0:0] pwr_vcore_ok,
    input [0:0] backup_protect,
// signals connected to CPU 
    input [0:0] c1_sleep,
    input [0:0] c2_sleep,
    input [0:0] c1_deepsleep,
    input [0:0] c2_deepsleep,
    output [0:0] rcc_c1_clk,
    output [0:0] rcc_c2_clk,
    output [0:0] rcc_fclk_c1,
    output [0:0] rcc_fclk_c2,
    output [0:0] rcc_c1_systick_clk,
    output [0:0] rcc_c2_systick_clk,
    output [0:0] rcc_c1_rst_n,
    output [0:0] rcc_c2_rst_n,
// signals connected to FLASH 
    output [0:0] rcc_obl_rst,
    output [0:0] rcc_obl_clk,
    output [0:0] rcc_flash_rst,
    output [0:0] rcc_flash_aclk,
    output [0:0] rcc_flash_hclk,
    input [0:0] flash_obl_reload,
    input [0:0] Tamp_rst_req,
    input [7:0] flash_csi_opt,
    input [11:0] flash_hsi_opt,
    input [0:0] obl_done,
// signals connected to CRS 
    input [9:0] crs_hsi48_trim,
// signals connected to 各类外设 
    output [0:0] rcc_perx_rst,
    output [0:0] rcc_perx_pclk,
    output [0:0] rcc_perx_hclk,
    output [0:0] rcc_perx_aclk,
    output [0:0] rcc_perx_ker_clk,
    input [0:0] perx_ker_clk_req,
// signals connected to 总线矩阵 
    output [0:0] rcc_axibridge_d1_clk,
    output [0:0] rcc_ahb3bridge_d1_clk,
    output [0:0] rcc_apb3bridge_d1_clk,
    output [0:0] rcc_ahb1bridge_d2_clk,
    output [0:0] rcc_ahb2bridge_d2_clk,
    output [0:0] rcc_apb1bridge_d2_clk,
    output [0:0] rcc_apb2bridge_d2_clk,
    output [0:0] rcc_ahb4bridge_d3_clk,
    output [0:0] rcc_apb4bridge_d3_clk,
    output [0:0] rcc_axibridge_rst,
    output [0:0] rcc_ahb3bridge_rst,
    output [0:0] rcc_apb3bridge_rst,
    output [0:0] rcc_ahb1bridge_rst,
    output [0:0] rcc_ahb2bridge_rst,
    output [0:0] rcc_apb1bridge_rst,
    output [0:0] rcc_apb2bridge_rst,
    output [0:0] rcc_ahb4bridge_rst,
    output [0:0] rcc_apb4bridge_rst,
    output [0:0] rcc_bus_clk_en,
// signals connected to 总线信号 
    input [0:0] RCCahblite总线信号,
// signals connected to 中断信号 
    output [0:0] rcc_it,
    output [0:0] rcc_hsecss_it,
    output [0:0] rcc_lsecss_it,
    output [0:0] rcc_hsecss_fail,
    output [0:0] rcc_lsecss_fail,
// signals connected to 复位源 
    input [0:0] iwdg1_out_rst,
    input [0:0] wwdg1_out_rst,
    input [0:0] iwdg2_out_rst,
    input [0:0] wwdg2_out_rst,
    input [0:0] lpwr1_rst,
    input [0:0] lpwr2_rst,
    input [0:0] pwr_bor_rst,
    input [0:0] pwr_por_rst,
    input [0:0] pwr_vsw_rst,
    input [0:0] d1_rst,
    input [0:0] d2_rst,
    input [0:0] stby_rst,
    input [0:0] cpu1_sftrst,
    input [0:0] cpu2_sftrst,
// signals connected to busy 指示信号 
    input [0:0] axibridge_d1_busy,
    input [0:0] ahbbridge_d1_busy,
    input [0:0] apbbridge_d1_busy,
    input [0:0] ahb1bridge_d2_busy,
    input [0:0] ahb2bridge_d2_busy,
    input [0:0] apb1bridge_d2_busy,
    input [0:0] apb2bridge_d2_busy,
    input [0:0] ahb4bridge_d3_busy,
    input [0:0] apb4bridge_d3_busy,
    input [0:0] flash_busy,
// signals connected to PLL * 3 
    input [0:0] pllx_rdy,
    output [0:0] pllx_on,
    output [0:0] divrx_en,
    output [0:0] divqx_en,
    output [0:0] divpx_en,
    output [1:0] pllx_rge,
    output [0:0] pllx_vco_sel,
    output [0:0] pllx_frac_en,
    output [6:0] rcc_pllx_divrx,
    output [6:0] rcc_pllx_divqx,
    output [6:0] rcc_pllx_divpx,
    output [8:0] rcc_pllx_divnx,
    output [12:0] rcc_pllx_fracnx,
    output [0:0] rcc_pllx_ref_clk,
    input [0:0] pllx_pclk,
    input [0:0] pllx_qclk,
    input [0:0] pllx_rclk,
// signals connected to HSE 
    output [0:0] hse_css_on,
    output [0:0] hse_byp,
    input [0:0] hse_rdy,
    output [0:0] hse_on,
    input [0:0] hse_css_fail,
    input [0:0] hse_clk,
// signals connected to HSI48 
    input [0:0] hsi48_ready,
    output [0:0] hsi48_on,
    output [9:0] hsi48_trim,
    input [0:0] hsi48_clk,
// signals connected to CSI 
    output [0:0] csi_on,
    input [0:0] csi_rdy,
    output [7:0] csi_trim,
    input [0:0] csi_clk,
// signals connected to HSI 
    input [0:0] hsi_rdy,
    output [0:0] hsi_on,
    output [11:0] hsi_trim,
    input [0:0] hsi_origin_clk,
// signals connected to LSE 
    input [0:0] lse_css_fail,
    output [0:0] lse_css_on,
    output [0:0] lse_drv,
    output [0:0] lse_byp,
    input [0:0] lse_rdy,
    output [0:0] lse_on,
    input [0:0] lse_clk,
// signals connected to LSI 
    input [0:0] lsi_rdy,
    output [0:0] lsi_on,
    input [0:0] lsi_clk,
);


 endmodule
